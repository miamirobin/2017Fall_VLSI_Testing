name bar
i a[0]
i a[1]
i a[2]
i a[3]
i a[4]
i a[5]
i a[6]
i a[7]
i a[8]
i a[9]
i a[10]
i a[11]
i a[12]
i a[13]
i a[14]
i a[15]
i a[16]
i a[17]
i a[18]
i a[19]
i a[20]
i a[21]
i a[22]
i a[23]
i a[24]
i a[25]
i a[26]
i a[27]
i a[28]
i a[29]
i a[30]
i a[31]
i a[32]
i a[33]
i a[34]
i a[35]
i a[36]
i a[37]
i a[38]
i a[39]
i a[40]
i a[41]
i a[42]
i a[43]
i a[44]
i a[45]
i a[46]
i a[47]
i a[48]
i a[49]
i a[50]
i a[51]
i a[52]
i a[53]
i a[54]
i a[55]
i a[56]
i a[57]
i a[58]
i a[59]
i a[60]
i a[61]
i a[62]
i a[63]
i a[64]
i a[65]
i a[66]
i a[67]
i a[68]
i a[69]
i a[70]
i a[71]
i a[72]
i a[73]
i a[74]
i a[75]
i a[76]
i a[77]
i a[78]
i a[79]
i a[80]
i a[81]
i a[82]
i a[83]
i a[84]
i a[85]
i a[86]
i a[87]
i a[88]
i a[89]
i a[90]
i a[91]
i a[92]
i a[93]
i a[94]
i a[95]
i a[96]
i a[97]
i a[98]
i a[99]
i a[100]
i a[101]
i a[102]
i a[103]
i a[104]
i a[105]
i a[106]
i a[107]
i a[108]
i a[109]
i a[110]
i a[111]
i a[112]
i a[113]
i a[114]
i a[115]
i a[116]
i a[117]
i a[118]
i a[119]
i a[120]
i a[121]
i a[122]
i a[123]
i a[124]
i a[125]
i a[126]
i a[127]
i shift[0]
i shift[1]
i shift[2]
i shift[3]
i shift[4]
i shift[5]
i shift[6]

g1 and a[77] shift[0] ; n264
g2 and shift[1] n264 ; n265
g3 and a[78] shift[0]_not ; n266
g4 and shift[1] n266 ; n267
g5 and n265_not n267_not ; n268
g6 and a[80] shift[0]_not ; n269
g7 and shift[1]_not n269 ; n270
g8 and a[79] shift[0] ; n271
g9 and shift[1]_not n271 ; n272
g10 and n270_not n272_not ; n273
g11 and n268 n273 ; n274
g12 and shift[2]_not shift[3]_not ; n275
g13 and n274_not n275 ; n276
g14 and a[73] shift[0] ; n277
g15 and shift[1] n277 ; n278
g16 and a[74] shift[0]_not ; n279
g17 and shift[1] n279 ; n280
g18 and n278_not n280_not ; n281
g19 and a[76] shift[0]_not ; n282
g20 and shift[1]_not n282 ; n283
g21 and a[75] shift[0] ; n284
g22 and shift[1]_not n284 ; n285
g23 and n283_not n285_not ; n286
g24 and n281 n286 ; n287
g25 and shift[2] shift[3]_not ; n288
g26 and n287_not n288 ; n289
g27 and n276_not n289_not ; n290
g28 and a[65] shift[0] ; n291
g29 and shift[1] n291 ; n292
g30 and a[66] shift[0]_not ; n293
g31 and shift[1] n293 ; n294
g32 and n292_not n294_not ; n295
g33 and a[68] shift[0]_not ; n296
g34 and shift[1]_not n296 ; n297
g35 and a[67] shift[0] ; n298
g36 and shift[1]_not n298 ; n299
g37 and n297_not n299_not ; n300
g38 and n295 n300 ; n301
g39 and shift[2] shift[3] ; n302
g40 and n301_not n302 ; n303
g41 and a[69] shift[0] ; n304
g42 and shift[1] n304 ; n305
g43 and a[70] shift[0]_not ; n306
g44 and shift[1] n306 ; n307
g45 and n305_not n307_not ; n308
g46 and a[72] shift[0]_not ; n309
g47 and shift[1]_not n309 ; n310
g48 and a[71] shift[0] ; n311
g49 and shift[1]_not n311 ; n312
g50 and n310_not n312_not ; n313
g51 and n308 n313 ; n314
g52 and shift[2]_not shift[3] ; n315
g53 and n314_not n315 ; n316
g54 and n303_not n316_not ; n317
g55 and n290 n317 ; n318
g56 and shift[4] shift[5] ; n319
g57 and n318_not n319 ; n320
g58 and a[93] shift[0] ; n321
g59 and shift[1] n321 ; n322
g60 and a[94] shift[0]_not ; n323
g61 and shift[1] n323 ; n324
g62 and n322_not n324_not ; n325
g63 and a[96] shift[0]_not ; n326
g64 and shift[1]_not n326 ; n327
g65 and a[95] shift[0] ; n328
g66 and shift[1]_not n328 ; n329
g67 and n327_not n329_not ; n330
g68 and n325 n330 ; n331
g69 and n275 n331_not ; n332
g70 and a[89] shift[0] ; n333
g71 and shift[1] n333 ; n334
g72 and a[90] shift[0]_not ; n335
g73 and shift[1] n335 ; n336
g74 and n334_not n336_not ; n337
g75 and a[92] shift[0]_not ; n338
g76 and shift[1]_not n338 ; n339
g77 and a[91] shift[0] ; n340
g78 and shift[1]_not n340 ; n341
g79 and n339_not n341_not ; n342
g80 and n337 n342 ; n343
g81 and n288 n343_not ; n344
g82 and n332_not n344_not ; n345
g83 and a[81] shift[0] ; n346
g84 and shift[1] n346 ; n347
g85 and a[82] shift[0]_not ; n348
g86 and shift[1] n348 ; n349
g87 and n347_not n349_not ; n350
g88 and a[84] shift[0]_not ; n351
g89 and shift[1]_not n351 ; n352
g90 and a[83] shift[0] ; n353
g91 and shift[1]_not n353 ; n354
g92 and n352_not n354_not ; n355
g93 and n350 n355 ; n356
g94 and n302 n356_not ; n357
g95 and a[85] shift[0] ; n358
g96 and shift[1] n358 ; n359
g97 and a[86] shift[0]_not ; n360
g98 and shift[1] n360 ; n361
g99 and n359_not n361_not ; n362
g100 and a[88] shift[0]_not ; n363
g101 and shift[1]_not n363 ; n364
g102 and a[87] shift[0] ; n365
g103 and shift[1]_not n365 ; n366
g104 and n364_not n366_not ; n367
g105 and n362 n367 ; n368
g106 and n315 n368_not ; n369
g107 and n357_not n369_not ; n370
g108 and n345 n370 ; n371
g109 and shift[4]_not shift[5] ; n372
g110 and n371_not n372 ; n373
g111 and n320_not n373_not ; n374
g112 and a[125] shift[0] ; n375
g113 and shift[1] n375 ; n376
g114 and a[126] shift[0]_not ; n377
g115 and shift[1] n377 ; n378
g116 and n376_not n378_not ; n379
g117 and a[0] shift[0]_not ; n380
g118 and shift[1]_not n380 ; n381
g119 and a[127] shift[0] ; n382
g120 and shift[1]_not n382 ; n383
g121 and n381_not n383_not ; n384
g122 and n379 n384 ; n385
g123 and n275 n385_not ; n386
g124 and a[121] shift[0] ; n387
g125 and shift[1] n387 ; n388
g126 and a[122] shift[0]_not ; n389
g127 and shift[1] n389 ; n390
g128 and n388_not n390_not ; n391
g129 and a[124] shift[0]_not ; n392
g130 and shift[1]_not n392 ; n393
g131 and a[123] shift[0] ; n394
g132 and shift[1]_not n394 ; n395
g133 and n393_not n395_not ; n396
g134 and n391 n396 ; n397
g135 and n288 n397_not ; n398
g136 and n386_not n398_not ; n399
g137 and a[113] shift[0] ; n400
g138 and shift[1] n400 ; n401
g139 and a[114] shift[0]_not ; n402
g140 and shift[1] n402 ; n403
g141 and n401_not n403_not ; n404
g142 and a[116] shift[0]_not ; n405
g143 and shift[1]_not n405 ; n406
g144 and a[115] shift[0] ; n407
g145 and shift[1]_not n407 ; n408
g146 and n406_not n408_not ; n409
g147 and n404 n409 ; n410
g148 and n302 n410_not ; n411
g149 and a[117] shift[0] ; n412
g150 and shift[1] n412 ; n413
g151 and a[118] shift[0]_not ; n414
g152 and shift[1] n414 ; n415
g153 and n413_not n415_not ; n416
g154 and a[120] shift[0]_not ; n417
g155 and shift[1]_not n417 ; n418
g156 and a[119] shift[0] ; n419
g157 and shift[1]_not n419 ; n420
g158 and n418_not n420_not ; n421
g159 and n416 n421 ; n422
g160 and n315 n422_not ; n423
g161 and n411_not n423_not ; n424
g162 and n399 n424 ; n425
g163 and shift[4]_not shift[5]_not ; n426
g164 and n425_not n426 ; n427
g165 and a[109] shift[0] ; n428
g166 and shift[1] n428 ; n429
g167 and a[110] shift[0]_not ; n430
g168 and shift[1] n430 ; n431
g169 and n429_not n431_not ; n432
g170 and a[112] shift[0]_not ; n433
g171 and shift[1]_not n433 ; n434
g172 and a[111] shift[0] ; n435
g173 and shift[1]_not n435 ; n436
g174 and n434_not n436_not ; n437
g175 and n432 n437 ; n438
g176 and n275 n438_not ; n439
g177 and a[105] shift[0] ; n440
g178 and shift[1] n440 ; n441
g179 and a[106] shift[0]_not ; n442
g180 and shift[1] n442 ; n443
g181 and n441_not n443_not ; n444
g182 and a[108] shift[0]_not ; n445
g183 and shift[1]_not n445 ; n446
g184 and a[107] shift[0] ; n447
g185 and shift[1]_not n447 ; n448
g186 and n446_not n448_not ; n449
g187 and n444 n449 ; n450
g188 and n288 n450_not ; n451
g189 and n439_not n451_not ; n452
g190 and a[97] shift[0] ; n453
g191 and shift[1] n453 ; n454
g192 and a[98] shift[0]_not ; n455
g193 and shift[1] n455 ; n456
g194 and n454_not n456_not ; n457
g195 and a[100] shift[0]_not ; n458
g196 and shift[1]_not n458 ; n459
g197 and a[99] shift[0] ; n460
g198 and shift[1]_not n460 ; n461
g199 and n459_not n461_not ; n462
g200 and n457 n462 ; n463
g201 and n302 n463_not ; n464
g202 and a[101] shift[0] ; n465
g203 and shift[1] n465 ; n466
g204 and a[102] shift[0]_not ; n467
g205 and shift[1] n467 ; n468
g206 and n466_not n468_not ; n469
g207 and a[104] shift[0]_not ; n470
g208 and shift[1]_not n470 ; n471
g209 and a[103] shift[0] ; n472
g210 and shift[1]_not n472 ; n473
g211 and n471_not n473_not ; n474
g212 and n469 n474 ; n475
g213 and n315 n475_not ; n476
g214 and n464_not n476_not ; n477
g215 and n452 n477 ; n478
g216 and shift[4] shift[5]_not ; n479
g217 and n478_not n479 ; n480
g218 and n427_not n480_not ; n481
g219 and n374 n481 ; n482
g220 and shift[6]_not n482_not ; n483
g221 and a[13] shift[0] ; n484
g222 and shift[1] n484 ; n485
g223 and a[14] shift[0]_not ; n486
g224 and shift[1] n486 ; n487
g225 and n485_not n487_not ; n488
g226 and a[16] shift[0]_not ; n489
g227 and shift[1]_not n489 ; n490
g228 and a[15] shift[0] ; n491
g229 and shift[1]_not n491 ; n492
g230 and n490_not n492_not ; n493
g231 and n488 n493 ; n494
g232 and n275 n494_not ; n495
g233 and a[9] shift[0] ; n496
g234 and shift[1] n496 ; n497
g235 and a[10] shift[0]_not ; n498
g236 and shift[1] n498 ; n499
g237 and n497_not n499_not ; n500
g238 and a[12] shift[0]_not ; n501
g239 and shift[1]_not n501 ; n502
g240 and a[11] shift[0] ; n503
g241 and shift[1]_not n503 ; n504
g242 and n502_not n504_not ; n505
g243 and n500 n505 ; n506
g244 and n288 n506_not ; n507
g245 and n495_not n507_not ; n508
g246 and a[1] shift[0] ; n509
g247 and shift[1] n509 ; n510
g248 and a[2] shift[0]_not ; n511
g249 and shift[1] n511 ; n512
g250 and n510_not n512_not ; n513
g251 and a[4] shift[0]_not ; n514
g252 and shift[1]_not n514 ; n515
g253 and a[3] shift[0] ; n516
g254 and shift[1]_not n516 ; n517
g255 and n515_not n517_not ; n518
g256 and n513 n518 ; n519
g257 and n302 n519_not ; n520
g258 and a[5] shift[0] ; n521
g259 and shift[1] n521 ; n522
g260 and a[6] shift[0]_not ; n523
g261 and shift[1] n523 ; n524
g262 and n522_not n524_not ; n525
g263 and a[8] shift[0]_not ; n526
g264 and shift[1]_not n526 ; n527
g265 and a[7] shift[0] ; n528
g266 and shift[1]_not n528 ; n529
g267 and n527_not n529_not ; n530
g268 and n525 n530 ; n531
g269 and n315 n531_not ; n532
g270 and n520_not n532_not ; n533
g271 and n508 n533 ; n534
g272 and n319 n534_not ; n535
g273 and a[29] shift[0] ; n536
g274 and shift[1] n536 ; n537
g275 and a[30] shift[0]_not ; n538
g276 and shift[1] n538 ; n539
g277 and n537_not n539_not ; n540
g278 and a[32] shift[0]_not ; n541
g279 and shift[1]_not n541 ; n542
g280 and a[31] shift[0] ; n543
g281 and shift[1]_not n543 ; n544
g282 and n542_not n544_not ; n545
g283 and n540 n545 ; n546
g284 and n275 n546_not ; n547
g285 and a[25] shift[0] ; n548
g286 and shift[1] n548 ; n549
g287 and a[26] shift[0]_not ; n550
g288 and shift[1] n550 ; n551
g289 and n549_not n551_not ; n552
g290 and a[28] shift[0]_not ; n553
g291 and shift[1]_not n553 ; n554
g292 and a[27] shift[0] ; n555
g293 and shift[1]_not n555 ; n556
g294 and n554_not n556_not ; n557
g295 and n552 n557 ; n558
g296 and n288 n558_not ; n559
g297 and n547_not n559_not ; n560
g298 and a[17] shift[0] ; n561
g299 and shift[1] n561 ; n562
g300 and a[18] shift[0]_not ; n563
g301 and shift[1] n563 ; n564
g302 and n562_not n564_not ; n565
g303 and a[20] shift[0]_not ; n566
g304 and shift[1]_not n566 ; n567
g305 and a[19] shift[0] ; n568
g306 and shift[1]_not n568 ; n569
g307 and n567_not n569_not ; n570
g308 and n565 n570 ; n571
g309 and n302 n571_not ; n572
g310 and a[21] shift[0] ; n573
g311 and shift[1] n573 ; n574
g312 and a[22] shift[0]_not ; n575
g313 and shift[1] n575 ; n576
g314 and n574_not n576_not ; n577
g315 and a[24] shift[0]_not ; n578
g316 and shift[1]_not n578 ; n579
g317 and a[23] shift[0] ; n580
g318 and shift[1]_not n580 ; n581
g319 and n579_not n581_not ; n582
g320 and n577 n582 ; n583
g321 and n315 n583_not ; n584
g322 and n572_not n584_not ; n585
g323 and n560 n585 ; n586
g324 and n372 n586_not ; n587
g325 and n535_not n587_not ; n588
g326 and a[61] shift[0] ; n589
g327 and shift[1] n589 ; n590
g328 and a[62] shift[0]_not ; n591
g329 and shift[1] n591 ; n592
g330 and n590_not n592_not ; n593
g331 and a[64] shift[0]_not ; n594
g332 and shift[1]_not n594 ; n595
g333 and a[63] shift[0] ; n596
g334 and shift[1]_not n596 ; n597
g335 and n595_not n597_not ; n598
g336 and n593 n598 ; n599
g337 and n275 n599_not ; n600
g338 and a[57] shift[0] ; n601
g339 and shift[1] n601 ; n602
g340 and a[58] shift[0]_not ; n603
g341 and shift[1] n603 ; n604
g342 and n602_not n604_not ; n605
g343 and a[60] shift[0]_not ; n606
g344 and shift[1]_not n606 ; n607
g345 and a[59] shift[0] ; n608
g346 and shift[1]_not n608 ; n609
g347 and n607_not n609_not ; n610
g348 and n605 n610 ; n611
g349 and n288 n611_not ; n612
g350 and n600_not n612_not ; n613
g351 and a[49] shift[0] ; n614
g352 and shift[1] n614 ; n615
g353 and a[50] shift[0]_not ; n616
g354 and shift[1] n616 ; n617
g355 and n615_not n617_not ; n618
g356 and a[52] shift[0]_not ; n619
g357 and shift[1]_not n619 ; n620
g358 and a[51] shift[0] ; n621
g359 and shift[1]_not n621 ; n622
g360 and n620_not n622_not ; n623
g361 and n618 n623 ; n624
g362 and n302 n624_not ; n625
g363 and a[53] shift[0] ; n626
g364 and shift[1] n626 ; n627
g365 and a[54] shift[0]_not ; n628
g366 and shift[1] n628 ; n629
g367 and n627_not n629_not ; n630
g368 and a[56] shift[0]_not ; n631
g369 and shift[1]_not n631 ; n632
g370 and a[55] shift[0] ; n633
g371 and shift[1]_not n633 ; n634
g372 and n632_not n634_not ; n635
g373 and n630 n635 ; n636
g374 and n315 n636_not ; n637
g375 and n625_not n637_not ; n638
g376 and n613 n638 ; n639
g377 and n426 n639_not ; n640
g378 and a[45] shift[0] ; n641
g379 and shift[1] n641 ; n642
g380 and a[46] shift[0]_not ; n643
g381 and shift[1] n643 ; n644
g382 and n642_not n644_not ; n645
g383 and a[48] shift[0]_not ; n646
g384 and shift[1]_not n646 ; n647
g385 and a[47] shift[0] ; n648
g386 and shift[1]_not n648 ; n649
g387 and n647_not n649_not ; n650
g388 and n645 n650 ; n651
g389 and n275 n651_not ; n652
g390 and a[41] shift[0] ; n653
g391 and shift[1] n653 ; n654
g392 and a[42] shift[0]_not ; n655
g393 and shift[1] n655 ; n656
g394 and n654_not n656_not ; n657
g395 and a[44] shift[0]_not ; n658
g396 and shift[1]_not n658 ; n659
g397 and a[43] shift[0] ; n660
g398 and shift[1]_not n660 ; n661
g399 and n659_not n661_not ; n662
g400 and n657 n662 ; n663
g401 and n288 n663_not ; n664
g402 and n652_not n664_not ; n665
g403 and a[33] shift[0] ; n666
g404 and shift[1] n666 ; n667
g405 and a[34] shift[0]_not ; n668
g406 and shift[1] n668 ; n669
g407 and n667_not n669_not ; n670
g408 and a[36] shift[0]_not ; n671
g409 and shift[1]_not n671 ; n672
g410 and a[35] shift[0] ; n673
g411 and shift[1]_not n673 ; n674
g412 and n672_not n674_not ; n675
g413 and n670 n675 ; n676
g414 and n302 n676_not ; n677
g415 and a[40] shift[0]_not ; n678
g416 and shift[1]_not n678 ; n679
g417 and a[37] shift[0] ; n680
g418 and shift[1] n680 ; n681
g419 and n679_not n681_not ; n682
g420 and a[39] shift[0] ; n683
g421 and shift[1]_not n683 ; n684
g422 and a[38] shift[0]_not ; n685
g423 and shift[1] n685 ; n686
g424 and n684_not n686_not ; n687
g425 and n682 n687 ; n688
g426 and n315 n688_not ; n689
g427 and n677_not n689_not ; n690
g428 and n665 n690 ; n691
g429 and n479 n691_not ; n692
g430 and n640_not n692_not ; n693
g431 and n588 n693 ; n694
g432 and shift[6] n694_not ; n695
g433 and n483_not n695_not ; result[0]
g434 and a[81] shift[0]_not ; n697
g435 and shift[1]_not n697 ; n698
g436 and a[78] shift[0] ; n699
g437 and shift[1] n699 ; n700
g438 and n698_not n700_not ; n701
g439 and a[80] shift[0] ; n702
g440 and shift[1]_not n702 ; n703
g441 and a[79] shift[0]_not ; n704
g442 and shift[1] n704 ; n705
g443 and n703_not n705_not ; n706
g444 and n701 n706 ; n707
g445 and n275 n707_not ; n708
g446 and a[77] shift[0]_not ; n709
g447 and shift[1]_not n709 ; n710
g448 and a[74] shift[0] ; n711
g449 and shift[1] n711 ; n712
g450 and n710_not n712_not ; n713
g451 and a[76] shift[0] ; n714
g452 and shift[1]_not n714 ; n715
g453 and a[75] shift[0]_not ; n716
g454 and shift[1] n716 ; n717
g455 and n715_not n717_not ; n718
g456 and n713 n718 ; n719
g457 and n288 n719_not ; n720
g458 and n708_not n720_not ; n721
g459 and a[69] shift[0]_not ; n722
g460 and shift[1]_not n722 ; n723
g461 and a[66] shift[0] ; n724
g462 and shift[1] n724 ; n725
g463 and n723_not n725_not ; n726
g464 and a[68] shift[0] ; n727
g465 and shift[1]_not n727 ; n728
g466 and a[67] shift[0]_not ; n729
g467 and shift[1] n729 ; n730
g468 and n728_not n730_not ; n731
g469 and n726 n731 ; n732
g470 and n302 n732_not ; n733
g471 and a[73] shift[0]_not ; n734
g472 and shift[1]_not n734 ; n735
g473 and a[70] shift[0] ; n736
g474 and shift[1] n736 ; n737
g475 and n735_not n737_not ; n738
g476 and a[72] shift[0] ; n739
g477 and shift[1]_not n739 ; n740
g478 and a[71] shift[0]_not ; n741
g479 and shift[1] n741 ; n742
g480 and n740_not n742_not ; n743
g481 and n738 n743 ; n744
g482 and n315 n744_not ; n745
g483 and n733_not n745_not ; n746
g484 and n721 n746 ; n747
g485 and n319 n747_not ; n748
g486 and a[97] shift[0]_not ; n749
g487 and shift[1]_not n749 ; n750
g488 and a[94] shift[0] ; n751
g489 and shift[1] n751 ; n752
g490 and n750_not n752_not ; n753
g491 and a[96] shift[0] ; n754
g492 and shift[1]_not n754 ; n755
g493 and a[95] shift[0]_not ; n756
g494 and shift[1] n756 ; n757
g495 and n755_not n757_not ; n758
g496 and n753 n758 ; n759
g497 and n275 n759_not ; n760
g498 and a[93] shift[0]_not ; n761
g499 and shift[1]_not n761 ; n762
g500 and a[90] shift[0] ; n763
g501 and shift[1] n763 ; n764
g502 and n762_not n764_not ; n765
g503 and a[92] shift[0] ; n766
g504 and shift[1]_not n766 ; n767
g505 and a[91] shift[0]_not ; n768
g506 and shift[1] n768 ; n769
g507 and n767_not n769_not ; n770
g508 and n765 n770 ; n771
g509 and n288 n771_not ; n772
g510 and n760_not n772_not ; n773
g511 and a[85] shift[0]_not ; n774
g512 and shift[1]_not n774 ; n775
g513 and a[82] shift[0] ; n776
g514 and shift[1] n776 ; n777
g515 and n775_not n777_not ; n778
g516 and a[84] shift[0] ; n779
g517 and shift[1]_not n779 ; n780
g518 and a[83] shift[0]_not ; n781
g519 and shift[1] n781 ; n782
g520 and n780_not n782_not ; n783
g521 and n778 n783 ; n784
g522 and n302 n784_not ; n785
g523 and a[89] shift[0]_not ; n786
g524 and shift[1]_not n786 ; n787
g525 and a[86] shift[0] ; n788
g526 and shift[1] n788 ; n789
g527 and n787_not n789_not ; n790
g528 and a[88] shift[0] ; n791
g529 and shift[1]_not n791 ; n792
g530 and a[87] shift[0]_not ; n793
g531 and shift[1] n793 ; n794
g532 and n792_not n794_not ; n795
g533 and n790 n795 ; n796
g534 and n315 n796_not ; n797
g535 and n785_not n797_not ; n798
g536 and n773 n798 ; n799
g537 and n372 n799_not ; n800
g538 and n748_not n800_not ; n801
g539 and a[1] shift[0]_not ; n802
g540 and shift[1]_not n802 ; n803
g541 and a[126] shift[0] ; n804
g542 and shift[1] n804 ; n805
g543 and n803_not n805_not ; n806
g544 and a[0] shift[0] ; n807
g545 and shift[1]_not n807 ; n808
g546 and a[127] shift[0]_not ; n809
g547 and shift[1] n809 ; n810
g548 and n808_not n810_not ; n811
g549 and n806 n811 ; n812
g550 and n275 n812_not ; n813
g551 and a[125] shift[0]_not ; n814
g552 and shift[1]_not n814 ; n815
g553 and a[122] shift[0] ; n816
g554 and shift[1] n816 ; n817
g555 and n815_not n817_not ; n818
g556 and a[124] shift[0] ; n819
g557 and shift[1]_not n819 ; n820
g558 and a[123] shift[0]_not ; n821
g559 and shift[1] n821 ; n822
g560 and n820_not n822_not ; n823
g561 and n818 n823 ; n824
g562 and n288 n824_not ; n825
g563 and n813_not n825_not ; n826
g564 and a[117] shift[0]_not ; n827
g565 and shift[1]_not n827 ; n828
g566 and a[114] shift[0] ; n829
g567 and shift[1] n829 ; n830
g568 and n828_not n830_not ; n831
g569 and a[116] shift[0] ; n832
g570 and shift[1]_not n832 ; n833
g571 and a[115] shift[0]_not ; n834
g572 and shift[1] n834 ; n835
g573 and n833_not n835_not ; n836
g574 and n831 n836 ; n837
g575 and n302 n837_not ; n838
g576 and a[121] shift[0]_not ; n839
g577 and shift[1]_not n839 ; n840
g578 and a[118] shift[0] ; n841
g579 and shift[1] n841 ; n842
g580 and n840_not n842_not ; n843
g581 and a[120] shift[0] ; n844
g582 and shift[1]_not n844 ; n845
g583 and a[119] shift[0]_not ; n846
g584 and shift[1] n846 ; n847
g585 and n845_not n847_not ; n848
g586 and n843 n848 ; n849
g587 and n315 n849_not ; n850
g588 and n838_not n850_not ; n851
g589 and n826 n851 ; n852
g590 and n426 n852_not ; n853
g591 and a[113] shift[0]_not ; n854
g592 and shift[1]_not n854 ; n855
g593 and a[110] shift[0] ; n856
g594 and shift[1] n856 ; n857
g595 and n855_not n857_not ; n858
g596 and a[112] shift[0] ; n859
g597 and shift[1]_not n859 ; n860
g598 and a[111] shift[0]_not ; n861
g599 and shift[1] n861 ; n862
g600 and n860_not n862_not ; n863
g601 and n858 n863 ; n864
g602 and n275 n864_not ; n865
g603 and a[109] shift[0]_not ; n866
g604 and shift[1]_not n866 ; n867
g605 and a[106] shift[0] ; n868
g606 and shift[1] n868 ; n869
g607 and n867_not n869_not ; n870
g608 and a[108] shift[0] ; n871
g609 and shift[1]_not n871 ; n872
g610 and a[107] shift[0]_not ; n873
g611 and shift[1] n873 ; n874
g612 and n872_not n874_not ; n875
g613 and n870 n875 ; n876
g614 and n288 n876_not ; n877
g615 and n865_not n877_not ; n878
g616 and a[101] shift[0]_not ; n879
g617 and shift[1]_not n879 ; n880
g618 and a[98] shift[0] ; n881
g619 and shift[1] n881 ; n882
g620 and n880_not n882_not ; n883
g621 and a[100] shift[0] ; n884
g622 and shift[1]_not n884 ; n885
g623 and a[99] shift[0]_not ; n886
g624 and shift[1] n886 ; n887
g625 and n885_not n887_not ; n888
g626 and n883 n888 ; n889
g627 and n302 n889_not ; n890
g628 and a[105] shift[0]_not ; n891
g629 and shift[1]_not n891 ; n892
g630 and a[102] shift[0] ; n893
g631 and shift[1] n893 ; n894
g632 and n892_not n894_not ; n895
g633 and a[104] shift[0] ; n896
g634 and shift[1]_not n896 ; n897
g635 and a[103] shift[0]_not ; n898
g636 and shift[1] n898 ; n899
g637 and n897_not n899_not ; n900
g638 and n895 n900 ; n901
g639 and n315 n901_not ; n902
g640 and n890_not n902_not ; n903
g641 and n878 n903 ; n904
g642 and n479 n904_not ; n905
g643 and n853_not n905_not ; n906
g644 and n801 n906 ; n907
g645 and shift[6]_not n907_not ; n908
g646 and a[65] shift[0]_not ; n909
g647 and shift[1]_not n909 ; n910
g648 and a[62] shift[0] ; n911
g649 and shift[1] n911 ; n912
g650 and n910_not n912_not ; n913
g651 and a[64] shift[0] ; n914
g652 and shift[1]_not n914 ; n915
g653 and a[63] shift[0]_not ; n916
g654 and shift[1] n916 ; n917
g655 and n915_not n917_not ; n918
g656 and n913 n918 ; n919
g657 and n275 n919_not ; n920
g658 and a[61] shift[0]_not ; n921
g659 and shift[1]_not n921 ; n922
g660 and a[58] shift[0] ; n923
g661 and shift[1] n923 ; n924
g662 and n922_not n924_not ; n925
g663 and a[60] shift[0] ; n926
g664 and shift[1]_not n926 ; n927
g665 and a[59] shift[0]_not ; n928
g666 and shift[1] n928 ; n929
g667 and n927_not n929_not ; n930
g668 and n925 n930 ; n931
g669 and n288 n931_not ; n932
g670 and n920_not n932_not ; n933
g671 and a[53] shift[0]_not ; n934
g672 and shift[1]_not n934 ; n935
g673 and a[50] shift[0] ; n936
g674 and shift[1] n936 ; n937
g675 and n935_not n937_not ; n938
g676 and a[52] shift[0] ; n939
g677 and shift[1]_not n939 ; n940
g678 and a[51] shift[0]_not ; n941
g679 and shift[1] n941 ; n942
g680 and n940_not n942_not ; n943
g681 and n938 n943 ; n944
g682 and n302 n944_not ; n945
g683 and a[57] shift[0]_not ; n946
g684 and shift[1]_not n946 ; n947
g685 and a[54] shift[0] ; n948
g686 and shift[1] n948 ; n949
g687 and n947_not n949_not ; n950
g688 and a[56] shift[0] ; n951
g689 and shift[1]_not n951 ; n952
g690 and a[55] shift[0]_not ; n953
g691 and shift[1] n953 ; n954
g692 and n952_not n954_not ; n955
g693 and n950 n955 ; n956
g694 and n315 n956_not ; n957
g695 and n945_not n957_not ; n958
g696 and n933 n958 ; n959
g697 and n426 n959_not ; n960
g698 and a[17] shift[0]_not ; n961
g699 and shift[1]_not n961 ; n962
g700 and a[14] shift[0] ; n963
g701 and shift[1] n963 ; n964
g702 and n962_not n964_not ; n965
g703 and a[16] shift[0] ; n966
g704 and shift[1]_not n966 ; n967
g705 and a[15] shift[0]_not ; n968
g706 and shift[1] n968 ; n969
g707 and n967_not n969_not ; n970
g708 and n965 n970 ; n971
g709 and n275 n971_not ; n972
g710 and a[13] shift[0]_not ; n973
g711 and shift[1]_not n973 ; n974
g712 and a[10] shift[0] ; n975
g713 and shift[1] n975 ; n976
g714 and n974_not n976_not ; n977
g715 and a[12] shift[0] ; n978
g716 and shift[1]_not n978 ; n979
g717 and a[11] shift[0]_not ; n980
g718 and shift[1] n980 ; n981
g719 and n979_not n981_not ; n982
g720 and n977 n982 ; n983
g721 and n288 n983_not ; n984
g722 and n972_not n984_not ; n985
g723 and a[5] shift[0]_not ; n986
g724 and shift[1]_not n986 ; n987
g725 and a[2] shift[0] ; n988
g726 and shift[1] n988 ; n989
g727 and n987_not n989_not ; n990
g728 and a[4] shift[0] ; n991
g729 and shift[1]_not n991 ; n992
g730 and a[3] shift[0]_not ; n993
g731 and shift[1] n993 ; n994
g732 and n992_not n994_not ; n995
g733 and n990 n995 ; n996
g734 and n302 n996_not ; n997
g735 and a[9] shift[0]_not ; n998
g736 and shift[1]_not n998 ; n999
g737 and a[6] shift[0] ; n1000
g738 and shift[1] n1000 ; n1001
g739 and n999_not n1001_not ; n1002
g740 and a[8] shift[0] ; n1003
g741 and shift[1]_not n1003 ; n1004
g742 and a[7] shift[0]_not ; n1005
g743 and shift[1] n1005 ; n1006
g744 and n1004_not n1006_not ; n1007
g745 and n1002 n1007 ; n1008
g746 and n315 n1008_not ; n1009
g747 and n997_not n1009_not ; n1010
g748 and n985 n1010 ; n1011
g749 and n319 n1011_not ; n1012
g750 and n960_not n1012_not ; n1013
g751 and a[49] shift[0]_not ; n1014
g752 and shift[1]_not n1014 ; n1015
g753 and a[46] shift[0] ; n1016
g754 and shift[1] n1016 ; n1017
g755 and n1015_not n1017_not ; n1018
g756 and a[48] shift[0] ; n1019
g757 and shift[1]_not n1019 ; n1020
g758 and a[47] shift[0]_not ; n1021
g759 and shift[1] n1021 ; n1022
g760 and n1020_not n1022_not ; n1023
g761 and n1018 n1023 ; n1024
g762 and n275 n1024_not ; n1025
g763 and a[42] shift[0] ; n1026
g764 and shift[1] n1026 ; n1027
g765 and a[43] shift[0]_not ; n1028
g766 and shift[1] n1028 ; n1029
g767 and n1027_not n1029_not ; n1030
g768 and a[45] shift[0]_not ; n1031
g769 and shift[1]_not n1031 ; n1032
g770 and a[44] shift[0] ; n1033
g771 and shift[1]_not n1033 ; n1034
g772 and n1032_not n1034_not ; n1035
g773 and n1030 n1035 ; n1036
g774 and n288 n1036_not ; n1037
g775 and n1025_not n1037_not ; n1038
g776 and a[37] shift[0]_not ; n1039
g777 and shift[1]_not n1039 ; n1040
g778 and a[34] shift[0] ; n1041
g779 and shift[1] n1041 ; n1042
g780 and n1040_not n1042_not ; n1043
g781 and a[36] shift[0] ; n1044
g782 and shift[1]_not n1044 ; n1045
g783 and a[35] shift[0]_not ; n1046
g784 and shift[1] n1046 ; n1047
g785 and n1045_not n1047_not ; n1048
g786 and n1043 n1048 ; n1049
g787 and n302 n1049_not ; n1050
g788 and a[41] shift[0]_not ; n1051
g789 and shift[1]_not n1051 ; n1052
g790 and a[40] shift[0] ; n1053
g791 and shift[1]_not n1053 ; n1054
g792 and n1052_not n1054_not ; n1055
g793 and a[39] shift[0]_not ; n1056
g794 and shift[1] n1056 ; n1057
g795 and a[38] shift[0] ; n1058
g796 and shift[1] n1058 ; n1059
g797 and n1057_not n1059_not ; n1060
g798 and n1055 n1060 ; n1061
g799 and n315 n1061_not ; n1062
g800 and n1050_not n1062_not ; n1063
g801 and n1038 n1063 ; n1064
g802 and n479 n1064_not ; n1065
g803 and a[33] shift[0]_not ; n1066
g804 and shift[1]_not n1066 ; n1067
g805 and a[30] shift[0] ; n1068
g806 and shift[1] n1068 ; n1069
g807 and n1067_not n1069_not ; n1070
g808 and a[32] shift[0] ; n1071
g809 and shift[1]_not n1071 ; n1072
g810 and a[31] shift[0]_not ; n1073
g811 and shift[1] n1073 ; n1074
g812 and n1072_not n1074_not ; n1075
g813 and n1070 n1075 ; n1076
g814 and n275 n1076_not ; n1077
g815 and a[29] shift[0]_not ; n1078
g816 and shift[1]_not n1078 ; n1079
g817 and a[26] shift[0] ; n1080
g818 and shift[1] n1080 ; n1081
g819 and n1079_not n1081_not ; n1082
g820 and a[28] shift[0] ; n1083
g821 and shift[1]_not n1083 ; n1084
g822 and a[27] shift[0]_not ; n1085
g823 and shift[1] n1085 ; n1086
g824 and n1084_not n1086_not ; n1087
g825 and n1082 n1087 ; n1088
g826 and n288 n1088_not ; n1089
g827 and n1077_not n1089_not ; n1090
g828 and a[21] shift[0]_not ; n1091
g829 and shift[1]_not n1091 ; n1092
g830 and a[18] shift[0] ; n1093
g831 and shift[1] n1093 ; n1094
g832 and n1092_not n1094_not ; n1095
g833 and a[20] shift[0] ; n1096
g834 and shift[1]_not n1096 ; n1097
g835 and a[19] shift[0]_not ; n1098
g836 and shift[1] n1098 ; n1099
g837 and n1097_not n1099_not ; n1100
g838 and n1095 n1100 ; n1101
g839 and n302 n1101_not ; n1102
g840 and a[25] shift[0]_not ; n1103
g841 and shift[1]_not n1103 ; n1104
g842 and a[22] shift[0] ; n1105
g843 and shift[1] n1105 ; n1106
g844 and n1104_not n1106_not ; n1107
g845 and a[24] shift[0] ; n1108
g846 and shift[1]_not n1108 ; n1109
g847 and a[23] shift[0]_not ; n1110
g848 and shift[1] n1110 ; n1111
g849 and n1109_not n1111_not ; n1112
g850 and n1107 n1112 ; n1113
g851 and n315 n1113_not ; n1114
g852 and n1102_not n1114_not ; n1115
g853 and n1090 n1115 ; n1116
g854 and n372 n1116_not ; n1117
g855 and n1065_not n1117_not ; n1118
g856 and n1013 n1118 ; n1119
g857 and shift[6] n1119_not ; n1120
g858 and n908_not n1120_not ; result[1]
g859 and shift[1]_not n346 ; n1122
g860 and shift[1]_not n348 ; n1123
g861 and n1122_not n1123_not ; n1124
g862 and shift[1] n269 ; n1125
g863 and shift[1] n271 ; n1126
g864 and n1125_not n1126_not ; n1127
g865 and n1124 n1127 ; n1128
g866 and n275 n1128_not ; n1129
g867 and shift[1]_not n264 ; n1130
g868 and shift[1]_not n266 ; n1131
g869 and n1130_not n1131_not ; n1132
g870 and shift[1] n282 ; n1133
g871 and shift[1] n284 ; n1134
g872 and n1133_not n1134_not ; n1135
g873 and n1132 n1135 ; n1136
g874 and n288 n1136_not ; n1137
g875 and n1129_not n1137_not ; n1138
g876 and shift[1]_not n304 ; n1139
g877 and shift[1]_not n306 ; n1140
g878 and n1139_not n1140_not ; n1141
g879 and shift[1] n296 ; n1142
g880 and shift[1] n298 ; n1143
g881 and n1142_not n1143_not ; n1144
g882 and n1141 n1144 ; n1145
g883 and n302 n1145_not ; n1146
g884 and shift[1]_not n277 ; n1147
g885 and shift[1]_not n279 ; n1148
g886 and n1147_not n1148_not ; n1149
g887 and shift[1] n309 ; n1150
g888 and shift[1] n311 ; n1151
g889 and n1150_not n1151_not ; n1152
g890 and n1149 n1152 ; n1153
g891 and n315 n1153_not ; n1154
g892 and n1146_not n1154_not ; n1155
g893 and n1138 n1155 ; n1156
g894 and n319 n1156_not ; n1157
g895 and shift[1]_not n453 ; n1158
g896 and shift[1]_not n455 ; n1159
g897 and n1158_not n1159_not ; n1160
g898 and shift[1] n326 ; n1161
g899 and shift[1] n328 ; n1162
g900 and n1161_not n1162_not ; n1163
g901 and n1160 n1163 ; n1164
g902 and n275 n1164_not ; n1165
g903 and shift[1]_not n321 ; n1166
g904 and shift[1]_not n323 ; n1167
g905 and n1166_not n1167_not ; n1168
g906 and shift[1] n338 ; n1169
g907 and shift[1] n340 ; n1170
g908 and n1169_not n1170_not ; n1171
g909 and n1168 n1171 ; n1172
g910 and n288 n1172_not ; n1173
g911 and n1165_not n1173_not ; n1174
g912 and shift[1]_not n358 ; n1175
g913 and shift[1]_not n360 ; n1176
g914 and n1175_not n1176_not ; n1177
g915 and shift[1] n351 ; n1178
g916 and shift[1] n353 ; n1179
g917 and n1178_not n1179_not ; n1180
g918 and n1177 n1180 ; n1181
g919 and n302 n1181_not ; n1182
g920 and shift[1]_not n333 ; n1183
g921 and shift[1]_not n335 ; n1184
g922 and n1183_not n1184_not ; n1185
g923 and shift[1] n363 ; n1186
g924 and shift[1] n365 ; n1187
g925 and n1186_not n1187_not ; n1188
g926 and n1185 n1188 ; n1189
g927 and n315 n1189_not ; n1190
g928 and n1182_not n1190_not ; n1191
g929 and n1174 n1191 ; n1192
g930 and n372 n1192_not ; n1193
g931 and n1157_not n1193_not ; n1194
g932 and shift[1]_not n509 ; n1195
g933 and shift[1]_not n511 ; n1196
g934 and n1195_not n1196_not ; n1197
g935 and shift[1] n380 ; n1198
g936 and shift[1] n382 ; n1199
g937 and n1198_not n1199_not ; n1200
g938 and n1197 n1200 ; n1201
g939 and n275 n1201_not ; n1202
g940 and shift[1]_not n375 ; n1203
g941 and shift[1]_not n377 ; n1204
g942 and n1203_not n1204_not ; n1205
g943 and shift[1] n392 ; n1206
g944 and shift[1] n394 ; n1207
g945 and n1206_not n1207_not ; n1208
g946 and n1205 n1208 ; n1209
g947 and n288 n1209_not ; n1210
g948 and n1202_not n1210_not ; n1211
g949 and shift[1]_not n412 ; n1212
g950 and shift[1]_not n414 ; n1213
g951 and n1212_not n1213_not ; n1214
g952 and shift[1] n405 ; n1215
g953 and shift[1] n407 ; n1216
g954 and n1215_not n1216_not ; n1217
g955 and n1214 n1217 ; n1218
g956 and n302 n1218_not ; n1219
g957 and shift[1]_not n387 ; n1220
g958 and shift[1]_not n389 ; n1221
g959 and n1220_not n1221_not ; n1222
g960 and shift[1] n417 ; n1223
g961 and shift[1] n419 ; n1224
g962 and n1223_not n1224_not ; n1225
g963 and n1222 n1225 ; n1226
g964 and n315 n1226_not ; n1227
g965 and n1219_not n1227_not ; n1228
g966 and n1211 n1228 ; n1229
g967 and n426 n1229_not ; n1230
g968 and shift[1]_not n400 ; n1231
g969 and shift[1]_not n402 ; n1232
g970 and n1231_not n1232_not ; n1233
g971 and shift[1] n433 ; n1234
g972 and shift[1] n435 ; n1235
g973 and n1234_not n1235_not ; n1236
g974 and n1233 n1236 ; n1237
g975 and n275 n1237_not ; n1238
g976 and shift[1]_not n428 ; n1239
g977 and shift[1]_not n430 ; n1240
g978 and n1239_not n1240_not ; n1241
g979 and shift[1] n445 ; n1242
g980 and shift[1] n447 ; n1243
g981 and n1242_not n1243_not ; n1244
g982 and n1241 n1244 ; n1245
g983 and n288 n1245_not ; n1246
g984 and n1238_not n1246_not ; n1247
g985 and shift[1]_not n465 ; n1248
g986 and shift[1]_not n467 ; n1249
g987 and n1248_not n1249_not ; n1250
g988 and shift[1] n458 ; n1251
g989 and shift[1] n460 ; n1252
g990 and n1251_not n1252_not ; n1253
g991 and n1250 n1253 ; n1254
g992 and n302 n1254_not ; n1255
g993 and shift[1]_not n440 ; n1256
g994 and shift[1]_not n442 ; n1257
g995 and n1256_not n1257_not ; n1258
g996 and shift[1] n470 ; n1259
g997 and shift[1] n472 ; n1260
g998 and n1259_not n1260_not ; n1261
g999 and n1258 n1261 ; n1262
g1000 and n315 n1262_not ; n1263
g1001 and n1255_not n1263_not ; n1264
g1002 and n1247 n1264 ; n1265
g1003 and n479 n1265_not ; n1266
g1004 and n1230_not n1266_not ; n1267
g1005 and n1194 n1267 ; n1268
g1006 and shift[6]_not n1268_not ; n1269
g1007 and shift[1]_not n291 ; n1270
g1008 and shift[1]_not n293 ; n1271
g1009 and n1270_not n1271_not ; n1272
g1010 and shift[1] n594 ; n1273
g1011 and shift[1] n596 ; n1274
g1012 and n1273_not n1274_not ; n1275
g1013 and n1272 n1275 ; n1276
g1014 and n275 n1276_not ; n1277
g1015 and shift[1]_not n589 ; n1278
g1016 and shift[1]_not n591 ; n1279
g1017 and n1278_not n1279_not ; n1280
g1018 and shift[1] n606 ; n1281
g1019 and shift[1] n608 ; n1282
g1020 and n1281_not n1282_not ; n1283
g1021 and n1280 n1283 ; n1284
g1022 and n288 n1284_not ; n1285
g1023 and n1277_not n1285_not ; n1286
g1024 and shift[1]_not n626 ; n1287
g1025 and shift[1]_not n628 ; n1288
g1026 and n1287_not n1288_not ; n1289
g1027 and shift[1] n619 ; n1290
g1028 and shift[1] n621 ; n1291
g1029 and n1290_not n1291_not ; n1292
g1030 and n1289 n1292 ; n1293
g1031 and n302 n1293_not ; n1294
g1032 and shift[1]_not n601 ; n1295
g1033 and shift[1]_not n603 ; n1296
g1034 and n1295_not n1296_not ; n1297
g1035 and shift[1] n631 ; n1298
g1036 and shift[1] n633 ; n1299
g1037 and n1298_not n1299_not ; n1300
g1038 and n1297 n1300 ; n1301
g1039 and n315 n1301_not ; n1302
g1040 and n1294_not n1302_not ; n1303
g1041 and n1286 n1303 ; n1304
g1042 and n426 n1304_not ; n1305
g1043 and shift[1]_not n561 ; n1306
g1044 and shift[1]_not n563 ; n1307
g1045 and n1306_not n1307_not ; n1308
g1046 and shift[1] n489 ; n1309
g1047 and shift[1] n491 ; n1310
g1048 and n1309_not n1310_not ; n1311
g1049 and n1308 n1311 ; n1312
g1050 and n275 n1312_not ; n1313
g1051 and shift[1]_not n484 ; n1314
g1052 and shift[1]_not n486 ; n1315
g1053 and n1314_not n1315_not ; n1316
g1054 and shift[1] n501 ; n1317
g1055 and shift[1] n503 ; n1318
g1056 and n1317_not n1318_not ; n1319
g1057 and n1316 n1319 ; n1320
g1058 and n288 n1320_not ; n1321
g1059 and n1313_not n1321_not ; n1322
g1060 and shift[1]_not n521 ; n1323
g1061 and shift[1]_not n523 ; n1324
g1062 and n1323_not n1324_not ; n1325
g1063 and shift[1] n514 ; n1326
g1064 and shift[1] n516 ; n1327
g1065 and n1326_not n1327_not ; n1328
g1066 and n1325 n1328 ; n1329
g1067 and n302 n1329_not ; n1330
g1068 and shift[1]_not n496 ; n1331
g1069 and shift[1]_not n498 ; n1332
g1070 and n1331_not n1332_not ; n1333
g1071 and shift[1] n526 ; n1334
g1072 and shift[1] n528 ; n1335
g1073 and n1334_not n1335_not ; n1336
g1074 and n1333 n1336 ; n1337
g1075 and n315 n1337_not ; n1338
g1076 and n1330_not n1338_not ; n1339
g1077 and n1322 n1339 ; n1340
g1078 and n319 n1340_not ; n1341
g1079 and n1305_not n1341_not ; n1342
g1080 and shift[1]_not n614 ; n1343
g1081 and shift[1]_not n616 ; n1344
g1082 and n1343_not n1344_not ; n1345
g1083 and shift[1] n646 ; n1346
g1084 and shift[1] n648 ; n1347
g1085 and n1346_not n1347_not ; n1348
g1086 and n1345 n1348 ; n1349
g1087 and n275 n1349_not ; n1350
g1088 and shift[1] n660 ; n1351
g1089 and shift[1] n658 ; n1352
g1090 and n1351_not n1352_not ; n1353
g1091 and shift[1]_not n643 ; n1354
g1092 and shift[1]_not n641 ; n1355
g1093 and n1354_not n1355_not ; n1356
g1094 and n1353 n1356 ; n1357
g1095 and n288 n1357_not ; n1358
g1096 and n1350_not n1358_not ; n1359
g1097 and shift[1]_not n680 ; n1360
g1098 and shift[1]_not n685 ; n1361
g1099 and n1360_not n1361_not ; n1362
g1100 and shift[1] n671 ; n1363
g1101 and shift[1] n673 ; n1364
g1102 and n1363_not n1364_not ; n1365
g1103 and n1362 n1365 ; n1366
g1104 and n302 n1366_not ; n1367
g1105 and shift[1]_not n653 ; n1368
g1106 and shift[1]_not n655 ; n1369
g1107 and n1368_not n1369_not ; n1370
g1108 and shift[1] n683 ; n1371
g1109 and shift[1] n678 ; n1372
g1110 and n1371_not n1372_not ; n1373
g1111 and n1370 n1373 ; n1374
g1112 and n315 n1374_not ; n1375
g1113 and n1367_not n1375_not ; n1376
g1114 and n1359 n1376 ; n1377
g1115 and n479 n1377_not ; n1378
g1116 and shift[1]_not n666 ; n1379
g1117 and shift[1]_not n668 ; n1380
g1118 and n1379_not n1380_not ; n1381
g1119 and shift[1] n541 ; n1382
g1120 and shift[1] n543 ; n1383
g1121 and n1382_not n1383_not ; n1384
g1122 and n1381 n1384 ; n1385
g1123 and n275 n1385_not ; n1386
g1124 and shift[1]_not n536 ; n1387
g1125 and shift[1]_not n538 ; n1388
g1126 and n1387_not n1388_not ; n1389
g1127 and shift[1] n553 ; n1390
g1128 and shift[1] n555 ; n1391
g1129 and n1390_not n1391_not ; n1392
g1130 and n1389 n1392 ; n1393
g1131 and n288 n1393_not ; n1394
g1132 and n1386_not n1394_not ; n1395
g1133 and shift[1]_not n573 ; n1396
g1134 and shift[1]_not n575 ; n1397
g1135 and n1396_not n1397_not ; n1398
g1136 and shift[1] n566 ; n1399
g1137 and shift[1] n568 ; n1400
g1138 and n1399_not n1400_not ; n1401
g1139 and n1398 n1401 ; n1402
g1140 and n302 n1402_not ; n1403
g1141 and shift[1]_not n548 ; n1404
g1142 and shift[1]_not n550 ; n1405
g1143 and n1404_not n1405_not ; n1406
g1144 and shift[1] n578 ; n1407
g1145 and shift[1] n580 ; n1408
g1146 and n1407_not n1408_not ; n1409
g1147 and n1406 n1409 ; n1410
g1148 and n315 n1410_not ; n1411
g1149 and n1403_not n1411_not ; n1412
g1150 and n1395 n1412 ; n1413
g1151 and n372 n1413_not ; n1414
g1152 and n1378_not n1414_not ; n1415
g1153 and n1342 n1415 ; n1416
g1154 and shift[6] n1416_not ; n1417
g1155 and n1269_not n1417_not ; result[2]
g1156 and shift[1] n854 ; n1419
g1157 and shift[1]_not n829 ; n1420
g1158 and n1419_not n1420_not ; n1421
g1159 and shift[1] n859 ; n1422
g1160 and shift[1]_not n834 ; n1423
g1161 and n1422_not n1423_not ; n1424
g1162 and n1421 n1424 ; n1425
g1163 and n275 n1425_not ; n1426
g1164 and shift[1] n866 ; n1427
g1165 and shift[1]_not n856 ; n1428
g1166 and n1427_not n1428_not ; n1429
g1167 and shift[1] n871 ; n1430
g1168 and shift[1]_not n861 ; n1431
g1169 and n1430_not n1431_not ; n1432
g1170 and n1429 n1432 ; n1433
g1171 and n288 n1433_not ; n1434
g1172 and n1426_not n1434_not ; n1435
g1173 and shift[1] n879 ; n1436
g1174 and shift[1]_not n893 ; n1437
g1175 and n1436_not n1437_not ; n1438
g1176 and shift[1] n884 ; n1439
g1177 and shift[1]_not n898 ; n1440
g1178 and n1439_not n1440_not ; n1441
g1179 and n1438 n1441 ; n1442
g1180 and n302 n1442_not ; n1443
g1181 and shift[1] n891 ; n1444
g1182 and shift[1]_not n868 ; n1445
g1183 and n1444_not n1445_not ; n1446
g1184 and shift[1] n896 ; n1447
g1185 and shift[1]_not n873 ; n1448
g1186 and n1447_not n1448_not ; n1449
g1187 and n1446 n1449 ; n1450
g1188 and n315 n1450_not ; n1451
g1189 and n1443_not n1451_not ; n1452
g1190 and n1435 n1452 ; n1453
g1191 and n479 n1453_not ; n1454
g1192 and shift[1] n749 ; n1455
g1193 and shift[1]_not n881 ; n1456
g1194 and n1455_not n1456_not ; n1457
g1195 and shift[1] n754 ; n1458
g1196 and shift[1]_not n886 ; n1459
g1197 and n1458_not n1459_not ; n1460
g1198 and n1457 n1460 ; n1461
g1199 and n275 n1461_not ; n1462
g1200 and shift[1] n761 ; n1463
g1201 and shift[1]_not n751 ; n1464
g1202 and n1463_not n1464_not ; n1465
g1203 and shift[1] n766 ; n1466
g1204 and shift[1]_not n756 ; n1467
g1205 and n1466_not n1467_not ; n1468
g1206 and n1465 n1468 ; n1469
g1207 and n288 n1469_not ; n1470
g1208 and n1462_not n1470_not ; n1471
g1209 and shift[1] n774 ; n1472
g1210 and shift[1]_not n788 ; n1473
g1211 and n1472_not n1473_not ; n1474
g1212 and shift[1] n779 ; n1475
g1213 and shift[1]_not n793 ; n1476
g1214 and n1475_not n1476_not ; n1477
g1215 and n1474 n1477 ; n1478
g1216 and n302 n1478_not ; n1479
g1217 and shift[1] n786 ; n1480
g1218 and shift[1]_not n763 ; n1481
g1219 and n1480_not n1481_not ; n1482
g1220 and shift[1] n791 ; n1483
g1221 and shift[1]_not n768 ; n1484
g1222 and n1483_not n1484_not ; n1485
g1223 and n1482 n1485 ; n1486
g1224 and n315 n1486_not ; n1487
g1225 and n1479_not n1487_not ; n1488
g1226 and n1471 n1488 ; n1489
g1227 and n372 n1489_not ; n1490
g1228 and n1454_not n1490_not ; n1491
g1229 and shift[1] n802 ; n1492
g1230 and shift[1]_not n988 ; n1493
g1231 and n1492_not n1493_not ; n1494
g1232 and shift[1] n807 ; n1495
g1233 and shift[1]_not n993 ; n1496
g1234 and n1495_not n1496_not ; n1497
g1235 and n1494 n1497 ; n1498
g1236 and n275 n1498_not ; n1499
g1237 and shift[1] n814 ; n1500
g1238 and shift[1]_not n804 ; n1501
g1239 and n1500_not n1501_not ; n1502
g1240 and shift[1] n819 ; n1503
g1241 and shift[1]_not n809 ; n1504
g1242 and n1503_not n1504_not ; n1505
g1243 and n1502 n1505 ; n1506
g1244 and n288 n1506_not ; n1507
g1245 and n1499_not n1507_not ; n1508
g1246 and shift[1] n827 ; n1509
g1247 and shift[1]_not n841 ; n1510
g1248 and n1509_not n1510_not ; n1511
g1249 and shift[1] n832 ; n1512
g1250 and shift[1]_not n846 ; n1513
g1251 and n1512_not n1513_not ; n1514
g1252 and n1511 n1514 ; n1515
g1253 and n302 n1515_not ; n1516
g1254 and shift[1] n839 ; n1517
g1255 and shift[1]_not n816 ; n1518
g1256 and n1517_not n1518_not ; n1519
g1257 and shift[1] n844 ; n1520
g1258 and shift[1]_not n821 ; n1521
g1259 and n1520_not n1521_not ; n1522
g1260 and n1519 n1522 ; n1523
g1261 and n315 n1523_not ; n1524
g1262 and n1516_not n1524_not ; n1525
g1263 and n1508 n1525 ; n1526
g1264 and n426 n1526_not ; n1527
g1265 and shift[1] n697 ; n1528
g1266 and shift[1]_not n776 ; n1529
g1267 and n1528_not n1529_not ; n1530
g1268 and shift[1] n702 ; n1531
g1269 and shift[1]_not n781 ; n1532
g1270 and n1531_not n1532_not ; n1533
g1271 and n1530 n1533 ; n1534
g1272 and n275 n1534_not ; n1535
g1273 and shift[1] n709 ; n1536
g1274 and shift[1]_not n699 ; n1537
g1275 and n1536_not n1537_not ; n1538
g1276 and shift[1] n714 ; n1539
g1277 and shift[1]_not n704 ; n1540
g1278 and n1539_not n1540_not ; n1541
g1279 and n1538 n1541 ; n1542
g1280 and n288 n1542_not ; n1543
g1281 and n1535_not n1543_not ; n1544
g1282 and shift[1] n722 ; n1545
g1283 and shift[1]_not n736 ; n1546
g1284 and n1545_not n1546_not ; n1547
g1285 and shift[1] n727 ; n1548
g1286 and shift[1]_not n741 ; n1549
g1287 and n1548_not n1549_not ; n1550
g1288 and n1547 n1550 ; n1551
g1289 and n302 n1551_not ; n1552
g1290 and shift[1] n734 ; n1553
g1291 and shift[1]_not n711 ; n1554
g1292 and n1553_not n1554_not ; n1555
g1293 and shift[1] n739 ; n1556
g1294 and shift[1]_not n716 ; n1557
g1295 and n1556_not n1557_not ; n1558
g1296 and n1555 n1558 ; n1559
g1297 and n315 n1559_not ; n1560
g1298 and n1552_not n1560_not ; n1561
g1299 and n1544 n1561 ; n1562
g1300 and n319 n1562_not ; n1563
g1301 and n1527_not n1563_not ; n1564
g1302 and n1491 n1564 ; n1565
g1303 and shift[6]_not n1565_not ; n1566
g1304 and shift[1] n909 ; n1567
g1305 and shift[1]_not n724 ; n1568
g1306 and n1567_not n1568_not ; n1569
g1307 and shift[1] n914 ; n1570
g1308 and shift[1]_not n729 ; n1571
g1309 and n1570_not n1571_not ; n1572
g1310 and n1569 n1572 ; n1573
g1311 and n275 n1573_not ; n1574
g1312 and shift[1] n921 ; n1575
g1313 and shift[1]_not n911 ; n1576
g1314 and n1575_not n1576_not ; n1577
g1315 and shift[1] n926 ; n1578
g1316 and shift[1]_not n916 ; n1579
g1317 and n1578_not n1579_not ; n1580
g1318 and n1577 n1580 ; n1581
g1319 and n288 n1581_not ; n1582
g1320 and n1574_not n1582_not ; n1583
g1321 and shift[1] n934 ; n1584
g1322 and shift[1]_not n948 ; n1585
g1323 and n1584_not n1585_not ; n1586
g1324 and shift[1] n939 ; n1587
g1325 and shift[1]_not n953 ; n1588
g1326 and n1587_not n1588_not ; n1589
g1327 and n1586 n1589 ; n1590
g1328 and n302 n1590_not ; n1591
g1329 and shift[1] n946 ; n1592
g1330 and shift[1]_not n923 ; n1593
g1331 and n1592_not n1593_not ; n1594
g1332 and shift[1] n951 ; n1595
g1333 and shift[1]_not n928 ; n1596
g1334 and n1595_not n1596_not ; n1597
g1335 and n1594 n1597 ; n1598
g1336 and n315 n1598_not ; n1599
g1337 and n1591_not n1599_not ; n1600
g1338 and n1583 n1600 ; n1601
g1339 and n426 n1601_not ; n1602
g1340 and shift[1] n1014 ; n1603
g1341 and shift[1]_not n936 ; n1604
g1342 and n1603_not n1604_not ; n1605
g1343 and shift[1] n1019 ; n1606
g1344 and shift[1]_not n941 ; n1607
g1345 and n1606_not n1607_not ; n1608
g1346 and n1605 n1608 ; n1609
g1347 and n275 n1609_not ; n1610
g1348 and shift[1] n1033 ; n1611
g1349 and shift[1] n1031 ; n1612
g1350 and n1611_not n1612_not ; n1613
g1351 and shift[1]_not n1021 ; n1614
g1352 and shift[1]_not n1016 ; n1615
g1353 and n1614_not n1615_not ; n1616
g1354 and n1613 n1616 ; n1617
g1355 and n288 n1617_not ; n1618
g1356 and n1610_not n1618_not ; n1619
g1357 and shift[1] n1039 ; n1620
g1358 and shift[1]_not n1058 ; n1621
g1359 and n1620_not n1621_not ; n1622
g1360 and shift[1] n1044 ; n1623
g1361 and shift[1]_not n1056 ; n1624
g1362 and n1623_not n1624_not ; n1625
g1363 and n1622 n1625 ; n1626
g1364 and n302 n1626_not ; n1627
g1365 and shift[1] n1051 ; n1628
g1366 and shift[1]_not n1026 ; n1629
g1367 and n1628_not n1629_not ; n1630
g1368 and shift[1] n1053 ; n1631
g1369 and shift[1]_not n1028 ; n1632
g1370 and n1631_not n1632_not ; n1633
g1371 and n1630 n1633 ; n1634
g1372 and n315 n1634_not ; n1635
g1373 and n1627_not n1635_not ; n1636
g1374 and n1619 n1636 ; n1637
g1375 and n479 n1637_not ; n1638
g1376 and n1602_not n1638_not ; n1639
g1377 and shift[1] n961 ; n1640
g1378 and shift[1]_not n1093 ; n1641
g1379 and n1640_not n1641_not ; n1642
g1380 and shift[1] n966 ; n1643
g1381 and shift[1]_not n1098 ; n1644
g1382 and n1643_not n1644_not ; n1645
g1383 and n1642 n1645 ; n1646
g1384 and n275 n1646_not ; n1647
g1385 and shift[1] n973 ; n1648
g1386 and shift[1]_not n963 ; n1649
g1387 and n1648_not n1649_not ; n1650
g1388 and shift[1] n978 ; n1651
g1389 and shift[1]_not n968 ; n1652
g1390 and n1651_not n1652_not ; n1653
g1391 and n1650 n1653 ; n1654
g1392 and n288 n1654_not ; n1655
g1393 and n1647_not n1655_not ; n1656
g1394 and shift[1] n986 ; n1657
g1395 and shift[1]_not n1000 ; n1658
g1396 and n1657_not n1658_not ; n1659
g1397 and shift[1] n991 ; n1660
g1398 and shift[1]_not n1005 ; n1661
g1399 and n1660_not n1661_not ; n1662
g1400 and n1659 n1662 ; n1663
g1401 and n302 n1663_not ; n1664
g1402 and shift[1] n998 ; n1665
g1403 and shift[1]_not n975 ; n1666
g1404 and n1665_not n1666_not ; n1667
g1405 and shift[1] n1003 ; n1668
g1406 and shift[1]_not n980 ; n1669
g1407 and n1668_not n1669_not ; n1670
g1408 and n1667 n1670 ; n1671
g1409 and n315 n1671_not ; n1672
g1410 and n1664_not n1672_not ; n1673
g1411 and n1656 n1673 ; n1674
g1412 and n319 n1674_not ; n1675
g1413 and shift[1] n1066 ; n1676
g1414 and shift[1]_not n1041 ; n1677
g1415 and n1676_not n1677_not ; n1678
g1416 and shift[1] n1071 ; n1679
g1417 and shift[1]_not n1046 ; n1680
g1418 and n1679_not n1680_not ; n1681
g1419 and n1678 n1681 ; n1682
g1420 and n275 n1682_not ; n1683
g1421 and shift[1] n1078 ; n1684
g1422 and shift[1]_not n1068 ; n1685
g1423 and n1684_not n1685_not ; n1686
g1424 and shift[1] n1083 ; n1687
g1425 and shift[1]_not n1073 ; n1688
g1426 and n1687_not n1688_not ; n1689
g1427 and n1686 n1689 ; n1690
g1428 and n288 n1690_not ; n1691
g1429 and n1683_not n1691_not ; n1692
g1430 and shift[1] n1091 ; n1693
g1431 and shift[1]_not n1105 ; n1694
g1432 and n1693_not n1694_not ; n1695
g1433 and shift[1] n1096 ; n1696
g1434 and shift[1]_not n1110 ; n1697
g1435 and n1696_not n1697_not ; n1698
g1436 and n1695 n1698 ; n1699
g1437 and n302 n1699_not ; n1700
g1438 and shift[1] n1103 ; n1701
g1439 and shift[1]_not n1080 ; n1702
g1440 and n1701_not n1702_not ; n1703
g1441 and shift[1] n1108 ; n1704
g1442 and shift[1]_not n1085 ; n1705
g1443 and n1704_not n1705_not ; n1706
g1444 and n1703 n1706 ; n1707
g1445 and n315 n1707_not ; n1708
g1446 and n1700_not n1708_not ; n1709
g1447 and n1692 n1709 ; n1710
g1448 and n372 n1710_not ; n1711
g1449 and n1675_not n1711_not ; n1712
g1450 and n1639 n1712 ; n1713
g1451 and shift[6] n1713_not ; n1714
g1452 and n1566_not n1714_not ; result[3]
g1453 and n275 n356_not ; n1716
g1454 and n274_not n288 ; n1717
g1455 and n1716_not n1717_not ; n1718
g1456 and n302 n314_not ; n1719
g1457 and n287_not n315 ; n1720
g1458 and n1719_not n1720_not ; n1721
g1459 and n1718 n1721 ; n1722
g1460 and n319 n1722_not ; n1723
g1461 and n275 n463_not ; n1724
g1462 and n288 n331_not ; n1725
g1463 and n1724_not n1725_not ; n1726
g1464 and n302 n368_not ; n1727
g1465 and n315 n343_not ; n1728
g1466 and n1727_not n1728_not ; n1729
g1467 and n1726 n1729 ; n1730
g1468 and n372 n1730_not ; n1731
g1469 and n1723_not n1731_not ; n1732
g1470 and n275 n519_not ; n1733
g1471 and n288 n385_not ; n1734
g1472 and n1733_not n1734_not ; n1735
g1473 and n302 n422_not ; n1736
g1474 and n315 n397_not ; n1737
g1475 and n1736_not n1737_not ; n1738
g1476 and n1735 n1738 ; n1739
g1477 and n426 n1739_not ; n1740
g1478 and n275 n410_not ; n1741
g1479 and n288 n438_not ; n1742
g1480 and n1741_not n1742_not ; n1743
g1481 and n302 n475_not ; n1744
g1482 and n315 n450_not ; n1745
g1483 and n1744_not n1745_not ; n1746
g1484 and n1743 n1746 ; n1747
g1485 and n479 n1747_not ; n1748
g1486 and n1740_not n1748_not ; n1749
g1487 and n1732 n1749 ; n1750
g1488 and shift[6]_not n1750_not ; n1751
g1489 and n275 n624_not ; n1752
g1490 and n288 n651_not ; n1753
g1491 and n1752_not n1753_not ; n1754
g1492 and n302 n688_not ; n1755
g1493 and n315 n663_not ; n1756
g1494 and n1755_not n1756_not ; n1757
g1495 and n1754 n1757 ; n1758
g1496 and n479 n1758_not ; n1759
g1497 and n275 n301_not ; n1760
g1498 and n288 n599_not ; n1761
g1499 and n1760_not n1761_not ; n1762
g1500 and n302 n636_not ; n1763
g1501 and n315 n611_not ; n1764
g1502 and n1763_not n1764_not ; n1765
g1503 and n1762 n1765 ; n1766
g1504 and n426 n1766_not ; n1767
g1505 and n1759_not n1767_not ; n1768
g1506 and n275 n676_not ; n1769
g1507 and n288 n546_not ; n1770
g1508 and n1769_not n1770_not ; n1771
g1509 and n302 n583_not ; n1772
g1510 and n315 n558_not ; n1773
g1511 and n1772_not n1773_not ; n1774
g1512 and n1771 n1774 ; n1775
g1513 and n372 n1775_not ; n1776
g1514 and n275 n571_not ; n1777
g1515 and n288 n494_not ; n1778
g1516 and n1777_not n1778_not ; n1779
g1517 and n302 n531_not ; n1780
g1518 and n315 n506_not ; n1781
g1519 and n1780_not n1781_not ; n1782
g1520 and n1779 n1782 ; n1783
g1521 and n319 n1783_not ; n1784
g1522 and n1776_not n1784_not ; n1785
g1523 and n1768 n1785 ; n1786
g1524 and shift[6] n1786_not ; n1787
g1525 and n1751_not n1787_not ; result[4]
g1526 and n275 n784_not ; n1789
g1527 and n288 n707_not ; n1790
g1528 and n1789_not n1790_not ; n1791
g1529 and n302 n744_not ; n1792
g1530 and n315 n719_not ; n1793
g1531 and n1792_not n1793_not ; n1794
g1532 and n1791 n1794 ; n1795
g1533 and n319 n1795_not ; n1796
g1534 and n275 n889_not ; n1797
g1535 and n288 n759_not ; n1798
g1536 and n1797_not n1798_not ; n1799
g1537 and n302 n796_not ; n1800
g1538 and n315 n771_not ; n1801
g1539 and n1800_not n1801_not ; n1802
g1540 and n1799 n1802 ; n1803
g1541 and n372 n1803_not ; n1804
g1542 and n1796_not n1804_not ; n1805
g1543 and n275 n996_not ; n1806
g1544 and n288 n812_not ; n1807
g1545 and n1806_not n1807_not ; n1808
g1546 and n302 n849_not ; n1809
g1547 and n315 n824_not ; n1810
g1548 and n1809_not n1810_not ; n1811
g1549 and n1808 n1811 ; n1812
g1550 and n426 n1812_not ; n1813
g1551 and n275 n837_not ; n1814
g1552 and n288 n864_not ; n1815
g1553 and n1814_not n1815_not ; n1816
g1554 and n302 n901_not ; n1817
g1555 and n315 n876_not ; n1818
g1556 and n1817_not n1818_not ; n1819
g1557 and n1816 n1819 ; n1820
g1558 and n479 n1820_not ; n1821
g1559 and n1813_not n1821_not ; n1822
g1560 and n1805 n1822 ; n1823
g1561 and shift[6]_not n1823_not ; n1824
g1562 and n275 n944_not ; n1825
g1563 and n288 n1024_not ; n1826
g1564 and n1825_not n1826_not ; n1827
g1565 and n302 n1061_not ; n1828
g1566 and n315 n1036_not ; n1829
g1567 and n1828_not n1829_not ; n1830
g1568 and n1827 n1830 ; n1831
g1569 and n479 n1831_not ; n1832
g1570 and n275 n732_not ; n1833
g1571 and n288 n919_not ; n1834
g1572 and n1833_not n1834_not ; n1835
g1573 and n302 n956_not ; n1836
g1574 and n315 n931_not ; n1837
g1575 and n1836_not n1837_not ; n1838
g1576 and n1835 n1838 ; n1839
g1577 and n426 n1839_not ; n1840
g1578 and n1832_not n1840_not ; n1841
g1579 and n275 n1049_not ; n1842
g1580 and n288 n1076_not ; n1843
g1581 and n1842_not n1843_not ; n1844
g1582 and n302 n1113_not ; n1845
g1583 and n315 n1088_not ; n1846
g1584 and n1845_not n1846_not ; n1847
g1585 and n1844 n1847 ; n1848
g1586 and n372 n1848_not ; n1849
g1587 and n275 n1101_not ; n1850
g1588 and n288 n971_not ; n1851
g1589 and n1850_not n1851_not ; n1852
g1590 and n302 n1008_not ; n1853
g1591 and n315 n983_not ; n1854
g1592 and n1853_not n1854_not ; n1855
g1593 and n1852 n1855 ; n1856
g1594 and n319 n1856_not ; n1857
g1595 and n1849_not n1857_not ; n1858
g1596 and n1841 n1858 ; n1859
g1597 and shift[6] n1859_not ; n1860
g1598 and n1824_not n1860_not ; result[5]
g1599 and n275 n1181_not ; n1862
g1600 and n288 n1128_not ; n1863
g1601 and n1862_not n1863_not ; n1864
g1602 and n302 n1153_not ; n1865
g1603 and n315 n1136_not ; n1866
g1604 and n1865_not n1866_not ; n1867
g1605 and n1864 n1867 ; n1868
g1606 and n319 n1868_not ; n1869
g1607 and n275 n1254_not ; n1870
g1608 and n288 n1164_not ; n1871
g1609 and n1870_not n1871_not ; n1872
g1610 and n302 n1189_not ; n1873
g1611 and n315 n1172_not ; n1874
g1612 and n1873_not n1874_not ; n1875
g1613 and n1872 n1875 ; n1876
g1614 and n372 n1876_not ; n1877
g1615 and n1869_not n1877_not ; n1878
g1616 and n275 n1329_not ; n1879
g1617 and n288 n1201_not ; n1880
g1618 and n1879_not n1880_not ; n1881
g1619 and n302 n1226_not ; n1882
g1620 and n315 n1209_not ; n1883
g1621 and n1882_not n1883_not ; n1884
g1622 and n1881 n1884 ; n1885
g1623 and n426 n1885_not ; n1886
g1624 and n275 n1218_not ; n1887
g1625 and n288 n1237_not ; n1888
g1626 and n1887_not n1888_not ; n1889
g1627 and n302 n1262_not ; n1890
g1628 and n315 n1245_not ; n1891
g1629 and n1890_not n1891_not ; n1892
g1630 and n1889 n1892 ; n1893
g1631 and n479 n1893_not ; n1894
g1632 and n1886_not n1894_not ; n1895
g1633 and n1878 n1895 ; n1896
g1634 and shift[6]_not n1896_not ; n1897
g1635 and n275 n1293_not ; n1898
g1636 and n288 n1349_not ; n1899
g1637 and n1898_not n1899_not ; n1900
g1638 and n302 n1374_not ; n1901
g1639 and n315 n1357_not ; n1902
g1640 and n1901_not n1902_not ; n1903
g1641 and n1900 n1903 ; n1904
g1642 and n479 n1904_not ; n1905
g1643 and n275 n1145_not ; n1906
g1644 and n288 n1276_not ; n1907
g1645 and n1906_not n1907_not ; n1908
g1646 and n302 n1301_not ; n1909
g1647 and n315 n1284_not ; n1910
g1648 and n1909_not n1910_not ; n1911
g1649 and n1908 n1911 ; n1912
g1650 and n426 n1912_not ; n1913
g1651 and n1905_not n1913_not ; n1914
g1652 and n275 n1366_not ; n1915
g1653 and n288 n1385_not ; n1916
g1654 and n1915_not n1916_not ; n1917
g1655 and n302 n1410_not ; n1918
g1656 and n315 n1393_not ; n1919
g1657 and n1918_not n1919_not ; n1920
g1658 and n1917 n1920 ; n1921
g1659 and n372 n1921_not ; n1922
g1660 and n275 n1402_not ; n1923
g1661 and n288 n1312_not ; n1924
g1662 and n1923_not n1924_not ; n1925
g1663 and n302 n1337_not ; n1926
g1664 and n315 n1320_not ; n1927
g1665 and n1926_not n1927_not ; n1928
g1666 and n1925 n1928 ; n1929
g1667 and n319 n1929_not ; n1930
g1668 and n1922_not n1930_not ; n1931
g1669 and n1914 n1931 ; n1932
g1670 and shift[6] n1932_not ; n1933
g1671 and n1897_not n1933_not ; result[6]
g1672 and n275 n1478_not ; n1935
g1673 and n288 n1534_not ; n1936
g1674 and n1935_not n1936_not ; n1937
g1675 and n302 n1559_not ; n1938
g1676 and n315 n1542_not ; n1939
g1677 and n1938_not n1939_not ; n1940
g1678 and n1937 n1940 ; n1941
g1679 and n319 n1941_not ; n1942
g1680 and n275 n1442_not ; n1943
g1681 and n288 n1461_not ; n1944
g1682 and n1943_not n1944_not ; n1945
g1683 and n302 n1486_not ; n1946
g1684 and n315 n1469_not ; n1947
g1685 and n1946_not n1947_not ; n1948
g1686 and n1945 n1948 ; n1949
g1687 and n372 n1949_not ; n1950
g1688 and n1942_not n1950_not ; n1951
g1689 and n275 n1663_not ; n1952
g1690 and n288 n1498_not ; n1953
g1691 and n1952_not n1953_not ; n1954
g1692 and n302 n1523_not ; n1955
g1693 and n315 n1506_not ; n1956
g1694 and n1955_not n1956_not ; n1957
g1695 and n1954 n1957 ; n1958
g1696 and n426 n1958_not ; n1959
g1697 and n275 n1515_not ; n1960
g1698 and n288 n1425_not ; n1961
g1699 and n1960_not n1961_not ; n1962
g1700 and n302 n1450_not ; n1963
g1701 and n315 n1433_not ; n1964
g1702 and n1963_not n1964_not ; n1965
g1703 and n1962 n1965 ; n1966
g1704 and n479 n1966_not ; n1967
g1705 and n1959_not n1967_not ; n1968
g1706 and n1951 n1968 ; n1969
g1707 and shift[6]_not n1969_not ; n1970
g1708 and n288 n1609_not ; n1971
g1709 and n315 n1617_not ; n1972
g1710 and n1971_not n1972_not ; n1973
g1711 and n302 n1634_not ; n1974
g1712 and n275 n1590_not ; n1975
g1713 and n1974_not n1975_not ; n1976
g1714 and n1973 n1976 ; n1977
g1715 and n479 n1977_not ; n1978
g1716 and n275 n1551_not ; n1979
g1717 and n288 n1573_not ; n1980
g1718 and n1979_not n1980_not ; n1981
g1719 and n302 n1598_not ; n1982
g1720 and n315 n1581_not ; n1983
g1721 and n1982_not n1983_not ; n1984
g1722 and n1981 n1984 ; n1985
g1723 and n426 n1985_not ; n1986
g1724 and n1978_not n1986_not ; n1987
g1725 and n275 n1626_not ; n1988
g1726 and n288 n1682_not ; n1989
g1727 and n1988_not n1989_not ; n1990
g1728 and n302 n1707_not ; n1991
g1729 and n315 n1690_not ; n1992
g1730 and n1991_not n1992_not ; n1993
g1731 and n1990 n1993 ; n1994
g1732 and n372 n1994_not ; n1995
g1733 and n275 n1699_not ; n1996
g1734 and n288 n1646_not ; n1997
g1735 and n1996_not n1997_not ; n1998
g1736 and n302 n1671_not ; n1999
g1737 and n315 n1654_not ; n2000
g1738 and n1999_not n2000_not ; n2001
g1739 and n1998 n2001 ; n2002
g1740 and n319 n2002_not ; n2003
g1741 and n1995_not n2003_not ; n2004
g1742 and n1987 n2004 ; n2005
g1743 and shift[6] n2005_not ; n2006
g1744 and n1970_not n2006_not ; result[7]
g1745 and n275 n368_not ; n2008
g1746 and n288 n356_not ; n2009
g1747 and n2008_not n2009_not ; n2010
g1748 and n287_not n302 ; n2011
g1749 and n274_not n315 ; n2012
g1750 and n2011_not n2012_not ; n2013
g1751 and n2010 n2013 ; n2014
g1752 and n319 n2014_not ; n2015
g1753 and n275 n475_not ; n2016
g1754 and n288 n463_not ; n2017
g1755 and n2016_not n2017_not ; n2018
g1756 and n302 n343_not ; n2019
g1757 and n315 n331_not ; n2020
g1758 and n2019_not n2020_not ; n2021
g1759 and n2018 n2021 ; n2022
g1760 and n372 n2022_not ; n2023
g1761 and n2015_not n2023_not ; n2024
g1762 and n275 n531_not ; n2025
g1763 and n288 n519_not ; n2026
g1764 and n2025_not n2026_not ; n2027
g1765 and n302 n397_not ; n2028
g1766 and n315 n385_not ; n2029
g1767 and n2028_not n2029_not ; n2030
g1768 and n2027 n2030 ; n2031
g1769 and n426 n2031_not ; n2032
g1770 and n275 n422_not ; n2033
g1771 and n288 n410_not ; n2034
g1772 and n2033_not n2034_not ; n2035
g1773 and n302 n450_not ; n2036
g1774 and n315 n438_not ; n2037
g1775 and n2036_not n2037_not ; n2038
g1776 and n2035 n2038 ; n2039
g1777 and n479 n2039_not ; n2040
g1778 and n2032_not n2040_not ; n2041
g1779 and n2024 n2041 ; n2042
g1780 and shift[6]_not n2042_not ; n2043
g1781 and n275 n636_not ; n2044
g1782 and n288 n624_not ; n2045
g1783 and n2044_not n2045_not ; n2046
g1784 and n302 n663_not ; n2047
g1785 and n315 n651_not ; n2048
g1786 and n2047_not n2048_not ; n2049
g1787 and n2046 n2049 ; n2050
g1788 and n479 n2050_not ; n2051
g1789 and n275 n314_not ; n2052
g1790 and n288 n301_not ; n2053
g1791 and n2052_not n2053_not ; n2054
g1792 and n302 n611_not ; n2055
g1793 and n315 n599_not ; n2056
g1794 and n2055_not n2056_not ; n2057
g1795 and n2054 n2057 ; n2058
g1796 and n426 n2058_not ; n2059
g1797 and n2051_not n2059_not ; n2060
g1798 and n275 n688_not ; n2061
g1799 and n288 n676_not ; n2062
g1800 and n2061_not n2062_not ; n2063
g1801 and n302 n558_not ; n2064
g1802 and n315 n546_not ; n2065
g1803 and n2064_not n2065_not ; n2066
g1804 and n2063 n2066 ; n2067
g1805 and n372 n2067_not ; n2068
g1806 and n275 n583_not ; n2069
g1807 and n288 n571_not ; n2070
g1808 and n2069_not n2070_not ; n2071
g1809 and n302 n506_not ; n2072
g1810 and n315 n494_not ; n2073
g1811 and n2072_not n2073_not ; n2074
g1812 and n2071 n2074 ; n2075
g1813 and n319 n2075_not ; n2076
g1814 and n2068_not n2076_not ; n2077
g1815 and n2060 n2077 ; n2078
g1816 and shift[6] n2078_not ; n2079
g1817 and n2043_not n2079_not ; result[8]
g1818 and n275 n796_not ; n2081
g1819 and n288 n784_not ; n2082
g1820 and n2081_not n2082_not ; n2083
g1821 and n302 n719_not ; n2084
g1822 and n315 n707_not ; n2085
g1823 and n2084_not n2085_not ; n2086
g1824 and n2083 n2086 ; n2087
g1825 and n319 n2087_not ; n2088
g1826 and n275 n901_not ; n2089
g1827 and n288 n889_not ; n2090
g1828 and n2089_not n2090_not ; n2091
g1829 and n302 n771_not ; n2092
g1830 and n315 n759_not ; n2093
g1831 and n2092_not n2093_not ; n2094
g1832 and n2091 n2094 ; n2095
g1833 and n372 n2095_not ; n2096
g1834 and n2088_not n2096_not ; n2097
g1835 and n275 n1008_not ; n2098
g1836 and n288 n996_not ; n2099
g1837 and n2098_not n2099_not ; n2100
g1838 and n302 n824_not ; n2101
g1839 and n315 n812_not ; n2102
g1840 and n2101_not n2102_not ; n2103
g1841 and n2100 n2103 ; n2104
g1842 and n426 n2104_not ; n2105
g1843 and n275 n849_not ; n2106
g1844 and n288 n837_not ; n2107
g1845 and n2106_not n2107_not ; n2108
g1846 and n302 n876_not ; n2109
g1847 and n315 n864_not ; n2110
g1848 and n2109_not n2110_not ; n2111
g1849 and n2108 n2111 ; n2112
g1850 and n479 n2112_not ; n2113
g1851 and n2105_not n2113_not ; n2114
g1852 and n2097 n2114 ; n2115
g1853 and shift[6]_not n2115_not ; n2116
g1854 and n275 n956_not ; n2117
g1855 and n288 n944_not ; n2118
g1856 and n2117_not n2118_not ; n2119
g1857 and n302 n1036_not ; n2120
g1858 and n315 n1024_not ; n2121
g1859 and n2120_not n2121_not ; n2122
g1860 and n2119 n2122 ; n2123
g1861 and n479 n2123_not ; n2124
g1862 and n275 n744_not ; n2125
g1863 and n288 n732_not ; n2126
g1864 and n2125_not n2126_not ; n2127
g1865 and n302 n931_not ; n2128
g1866 and n315 n919_not ; n2129
g1867 and n2128_not n2129_not ; n2130
g1868 and n2127 n2130 ; n2131
g1869 and n426 n2131_not ; n2132
g1870 and n2124_not n2132_not ; n2133
g1871 and n275 n1061_not ; n2134
g1872 and n288 n1049_not ; n2135
g1873 and n2134_not n2135_not ; n2136
g1874 and n302 n1088_not ; n2137
g1875 and n315 n1076_not ; n2138
g1876 and n2137_not n2138_not ; n2139
g1877 and n2136 n2139 ; n2140
g1878 and n372 n2140_not ; n2141
g1879 and n275 n1113_not ; n2142
g1880 and n288 n1101_not ; n2143
g1881 and n2142_not n2143_not ; n2144
g1882 and n302 n983_not ; n2145
g1883 and n315 n971_not ; n2146
g1884 and n2145_not n2146_not ; n2147
g1885 and n2144 n2147 ; n2148
g1886 and n319 n2148_not ; n2149
g1887 and n2141_not n2149_not ; n2150
g1888 and n2133 n2150 ; n2151
g1889 and shift[6] n2151_not ; n2152
g1890 and n2116_not n2152_not ; result[9]
g1891 and n275 n1189_not ; n2154
g1892 and n288 n1181_not ; n2155
g1893 and n2154_not n2155_not ; n2156
g1894 and n302 n1136_not ; n2157
g1895 and n315 n1128_not ; n2158
g1896 and n2157_not n2158_not ; n2159
g1897 and n2156 n2159 ; n2160
g1898 and n319 n2160_not ; n2161
g1899 and n275 n1262_not ; n2162
g1900 and n288 n1254_not ; n2163
g1901 and n2162_not n2163_not ; n2164
g1902 and n302 n1172_not ; n2165
g1903 and n315 n1164_not ; n2166
g1904 and n2165_not n2166_not ; n2167
g1905 and n2164 n2167 ; n2168
g1906 and n372 n2168_not ; n2169
g1907 and n2161_not n2169_not ; n2170
g1908 and n275 n1337_not ; n2171
g1909 and n288 n1329_not ; n2172
g1910 and n2171_not n2172_not ; n2173
g1911 and n302 n1209_not ; n2174
g1912 and n315 n1201_not ; n2175
g1913 and n2174_not n2175_not ; n2176
g1914 and n2173 n2176 ; n2177
g1915 and n426 n2177_not ; n2178
g1916 and n275 n1226_not ; n2179
g1917 and n288 n1218_not ; n2180
g1918 and n2179_not n2180_not ; n2181
g1919 and n302 n1245_not ; n2182
g1920 and n315 n1237_not ; n2183
g1921 and n2182_not n2183_not ; n2184
g1922 and n2181 n2184 ; n2185
g1923 and n479 n2185_not ; n2186
g1924 and n2178_not n2186_not ; n2187
g1925 and n2170 n2187 ; n2188
g1926 and shift[6]_not n2188_not ; n2189
g1927 and n275 n1301_not ; n2190
g1928 and n288 n1293_not ; n2191
g1929 and n2190_not n2191_not ; n2192
g1930 and n302 n1357_not ; n2193
g1931 and n315 n1349_not ; n2194
g1932 and n2193_not n2194_not ; n2195
g1933 and n2192 n2195 ; n2196
g1934 and n479 n2196_not ; n2197
g1935 and n275 n1153_not ; n2198
g1936 and n288 n1145_not ; n2199
g1937 and n2198_not n2199_not ; n2200
g1938 and n302 n1284_not ; n2201
g1939 and n315 n1276_not ; n2202
g1940 and n2201_not n2202_not ; n2203
g1941 and n2200 n2203 ; n2204
g1942 and n426 n2204_not ; n2205
g1943 and n2197_not n2205_not ; n2206
g1944 and n275 n1374_not ; n2207
g1945 and n288 n1366_not ; n2208
g1946 and n2207_not n2208_not ; n2209
g1947 and n302 n1393_not ; n2210
g1948 and n315 n1385_not ; n2211
g1949 and n2210_not n2211_not ; n2212
g1950 and n2209 n2212 ; n2213
g1951 and n372 n2213_not ; n2214
g1952 and n275 n1410_not ; n2215
g1953 and n288 n1402_not ; n2216
g1954 and n2215_not n2216_not ; n2217
g1955 and n302 n1320_not ; n2218
g1956 and n315 n1312_not ; n2219
g1957 and n2218_not n2219_not ; n2220
g1958 and n2217 n2220 ; n2221
g1959 and n319 n2221_not ; n2222
g1960 and n2214_not n2222_not ; n2223
g1961 and n2206 n2223 ; n2224
g1962 and shift[6] n2224_not ; n2225
g1963 and n2189_not n2225_not ; result[10]
g1964 and n275 n1486_not ; n2227
g1965 and n288 n1478_not ; n2228
g1966 and n2227_not n2228_not ; n2229
g1967 and n302 n1542_not ; n2230
g1968 and n315 n1534_not ; n2231
g1969 and n2230_not n2231_not ; n2232
g1970 and n2229 n2232 ; n2233
g1971 and n319 n2233_not ; n2234
g1972 and n275 n1450_not ; n2235
g1973 and n288 n1442_not ; n2236
g1974 and n2235_not n2236_not ; n2237
g1975 and n302 n1469_not ; n2238
g1976 and n315 n1461_not ; n2239
g1977 and n2238_not n2239_not ; n2240
g1978 and n2237 n2240 ; n2241
g1979 and n372 n2241_not ; n2242
g1980 and n2234_not n2242_not ; n2243
g1981 and n275 n1671_not ; n2244
g1982 and n288 n1663_not ; n2245
g1983 and n2244_not n2245_not ; n2246
g1984 and n302 n1506_not ; n2247
g1985 and n315 n1498_not ; n2248
g1986 and n2247_not n2248_not ; n2249
g1987 and n2246 n2249 ; n2250
g1988 and n426 n2250_not ; n2251
g1989 and n275 n1523_not ; n2252
g1990 and n288 n1515_not ; n2253
g1991 and n2252_not n2253_not ; n2254
g1992 and n302 n1433_not ; n2255
g1993 and n315 n1425_not ; n2256
g1994 and n2255_not n2256_not ; n2257
g1995 and n2254 n2257 ; n2258
g1996 and n479 n2258_not ; n2259
g1997 and n2251_not n2259_not ; n2260
g1998 and n2243 n2260 ; n2261
g1999 and shift[6]_not n2261_not ; n2262
g2000 and n275 n1598_not ; n2263
g2001 and n315 n1609_not ; n2264
g2002 and n2263_not n2264_not ; n2265
g2003 and n302 n1617_not ; n2266
g2004 and n288 n1590_not ; n2267
g2005 and n2266_not n2267_not ; n2268
g2006 and n2265 n2268 ; n2269
g2007 and n479 n2269_not ; n2270
g2008 and n275 n1559_not ; n2271
g2009 and n288 n1551_not ; n2272
g2010 and n2271_not n2272_not ; n2273
g2011 and n302 n1581_not ; n2274
g2012 and n315 n1573_not ; n2275
g2013 and n2274_not n2275_not ; n2276
g2014 and n2273 n2276 ; n2277
g2015 and n426 n2277_not ; n2278
g2016 and n2270_not n2278_not ; n2279
g2017 and n275 n1634_not ; n2280
g2018 and n288 n1626_not ; n2281
g2019 and n2280_not n2281_not ; n2282
g2020 and n302 n1690_not ; n2283
g2021 and n315 n1682_not ; n2284
g2022 and n2283_not n2284_not ; n2285
g2023 and n2282 n2285 ; n2286
g2024 and n372 n2286_not ; n2287
g2025 and n275 n1707_not ; n2288
g2026 and n288 n1699_not ; n2289
g2027 and n2288_not n2289_not ; n2290
g2028 and n302 n1654_not ; n2291
g2029 and n315 n1646_not ; n2292
g2030 and n2291_not n2292_not ; n2293
g2031 and n2290 n2293 ; n2294
g2032 and n319 n2294_not ; n2295
g2033 and n2287_not n2295_not ; n2296
g2034 and n2279 n2296 ; n2297
g2035 and shift[6] n2297_not ; n2298
g2036 and n2262_not n2298_not ; result[11]
g2037 and n275 n343_not ; n2300
g2038 and n288 n368_not ; n2301
g2039 and n2300_not n2301_not ; n2302
g2040 and n274_not n302 ; n2303
g2041 and n315 n356_not ; n2304
g2042 and n2303_not n2304_not ; n2305
g2043 and n2302 n2305 ; n2306
g2044 and n319 n2306_not ; n2307
g2045 and n275 n450_not ; n2308
g2046 and n288 n475_not ; n2309
g2047 and n2308_not n2309_not ; n2310
g2048 and n302 n331_not ; n2311
g2049 and n315 n463_not ; n2312
g2050 and n2311_not n2312_not ; n2313
g2051 and n2310 n2313 ; n2314
g2052 and n372 n2314_not ; n2315
g2053 and n2307_not n2315_not ; n2316
g2054 and n275 n506_not ; n2317
g2055 and n288 n531_not ; n2318
g2056 and n2317_not n2318_not ; n2319
g2057 and n302 n385_not ; n2320
g2058 and n315 n519_not ; n2321
g2059 and n2320_not n2321_not ; n2322
g2060 and n2319 n2322 ; n2323
g2061 and n426 n2323_not ; n2324
g2062 and n275 n397_not ; n2325
g2063 and n288 n422_not ; n2326
g2064 and n2325_not n2326_not ; n2327
g2065 and n302 n438_not ; n2328
g2066 and n315 n410_not ; n2329
g2067 and n2328_not n2329_not ; n2330
g2068 and n2327 n2330 ; n2331
g2069 and n479 n2331_not ; n2332
g2070 and n2324_not n2332_not ; n2333
g2071 and n2316 n2333 ; n2334
g2072 and shift[6]_not n2334_not ; n2335
g2073 and n275 n611_not ; n2336
g2074 and n288 n636_not ; n2337
g2075 and n2336_not n2337_not ; n2338
g2076 and n302 n651_not ; n2339
g2077 and n315 n624_not ; n2340
g2078 and n2339_not n2340_not ; n2341
g2079 and n2338 n2341 ; n2342
g2080 and n479 n2342_not ; n2343
g2081 and n275 n287_not ; n2344
g2082 and n288 n314_not ; n2345
g2083 and n2344_not n2345_not ; n2346
g2084 and n302 n599_not ; n2347
g2085 and n301_not n315 ; n2348
g2086 and n2347_not n2348_not ; n2349
g2087 and n2346 n2349 ; n2350
g2088 and n426 n2350_not ; n2351
g2089 and n2343_not n2351_not ; n2352
g2090 and n275 n663_not ; n2353
g2091 and n288 n688_not ; n2354
g2092 and n2353_not n2354_not ; n2355
g2093 and n302 n546_not ; n2356
g2094 and n315 n676_not ; n2357
g2095 and n2356_not n2357_not ; n2358
g2096 and n2355 n2358 ; n2359
g2097 and n372 n2359_not ; n2360
g2098 and n275 n558_not ; n2361
g2099 and n288 n583_not ; n2362
g2100 and n2361_not n2362_not ; n2363
g2101 and n302 n494_not ; n2364
g2102 and n315 n571_not ; n2365
g2103 and n2364_not n2365_not ; n2366
g2104 and n2363 n2366 ; n2367
g2105 and n319 n2367_not ; n2368
g2106 and n2360_not n2368_not ; n2369
g2107 and n2352 n2369 ; n2370
g2108 and shift[6] n2370_not ; n2371
g2109 and n2335_not n2371_not ; result[12]
g2110 and n275 n771_not ; n2373
g2111 and n288 n796_not ; n2374
g2112 and n2373_not n2374_not ; n2375
g2113 and n302 n707_not ; n2376
g2114 and n315 n784_not ; n2377
g2115 and n2376_not n2377_not ; n2378
g2116 and n2375 n2378 ; n2379
g2117 and n319 n2379_not ; n2380
g2118 and n275 n876_not ; n2381
g2119 and n288 n901_not ; n2382
g2120 and n2381_not n2382_not ; n2383
g2121 and n302 n759_not ; n2384
g2122 and n315 n889_not ; n2385
g2123 and n2384_not n2385_not ; n2386
g2124 and n2383 n2386 ; n2387
g2125 and n372 n2387_not ; n2388
g2126 and n2380_not n2388_not ; n2389
g2127 and n275 n983_not ; n2390
g2128 and n288 n1008_not ; n2391
g2129 and n2390_not n2391_not ; n2392
g2130 and n302 n812_not ; n2393
g2131 and n315 n996_not ; n2394
g2132 and n2393_not n2394_not ; n2395
g2133 and n2392 n2395 ; n2396
g2134 and n426 n2396_not ; n2397
g2135 and n275 n824_not ; n2398
g2136 and n288 n849_not ; n2399
g2137 and n2398_not n2399_not ; n2400
g2138 and n302 n864_not ; n2401
g2139 and n315 n837_not ; n2402
g2140 and n2401_not n2402_not ; n2403
g2141 and n2400 n2403 ; n2404
g2142 and n479 n2404_not ; n2405
g2143 and n2397_not n2405_not ; n2406
g2144 and n2389 n2406 ; n2407
g2145 and shift[6]_not n2407_not ; n2408
g2146 and n275 n931_not ; n2409
g2147 and n288 n956_not ; n2410
g2148 and n2409_not n2410_not ; n2411
g2149 and n302 n1024_not ; n2412
g2150 and n315 n944_not ; n2413
g2151 and n2412_not n2413_not ; n2414
g2152 and n2411 n2414 ; n2415
g2153 and n479 n2415_not ; n2416
g2154 and n275 n719_not ; n2417
g2155 and n288 n744_not ; n2418
g2156 and n2417_not n2418_not ; n2419
g2157 and n302 n919_not ; n2420
g2158 and n315 n732_not ; n2421
g2159 and n2420_not n2421_not ; n2422
g2160 and n2419 n2422 ; n2423
g2161 and n426 n2423_not ; n2424
g2162 and n2416_not n2424_not ; n2425
g2163 and n275 n1036_not ; n2426
g2164 and n288 n1061_not ; n2427
g2165 and n2426_not n2427_not ; n2428
g2166 and n302 n1076_not ; n2429
g2167 and n315 n1049_not ; n2430
g2168 and n2429_not n2430_not ; n2431
g2169 and n2428 n2431 ; n2432
g2170 and n372 n2432_not ; n2433
g2171 and n275 n1088_not ; n2434
g2172 and n288 n1113_not ; n2435
g2173 and n2434_not n2435_not ; n2436
g2174 and n302 n971_not ; n2437
g2175 and n315 n1101_not ; n2438
g2176 and n2437_not n2438_not ; n2439
g2177 and n2436 n2439 ; n2440
g2178 and n319 n2440_not ; n2441
g2179 and n2433_not n2441_not ; n2442
g2180 and n2425 n2442 ; n2443
g2181 and shift[6] n2443_not ; n2444
g2182 and n2408_not n2444_not ; result[13]
g2183 and n275 n1172_not ; n2446
g2184 and n288 n1189_not ; n2447
g2185 and n2446_not n2447_not ; n2448
g2186 and n302 n1128_not ; n2449
g2187 and n315 n1181_not ; n2450
g2188 and n2449_not n2450_not ; n2451
g2189 and n2448 n2451 ; n2452
g2190 and n319 n2452_not ; n2453
g2191 and n275 n1245_not ; n2454
g2192 and n288 n1262_not ; n2455
g2193 and n2454_not n2455_not ; n2456
g2194 and n302 n1164_not ; n2457
g2195 and n315 n1254_not ; n2458
g2196 and n2457_not n2458_not ; n2459
g2197 and n2456 n2459 ; n2460
g2198 and n372 n2460_not ; n2461
g2199 and n2453_not n2461_not ; n2462
g2200 and n275 n1320_not ; n2463
g2201 and n288 n1337_not ; n2464
g2202 and n2463_not n2464_not ; n2465
g2203 and n302 n1201_not ; n2466
g2204 and n315 n1329_not ; n2467
g2205 and n2466_not n2467_not ; n2468
g2206 and n2465 n2468 ; n2469
g2207 and n426 n2469_not ; n2470
g2208 and n275 n1209_not ; n2471
g2209 and n288 n1226_not ; n2472
g2210 and n2471_not n2472_not ; n2473
g2211 and n302 n1237_not ; n2474
g2212 and n315 n1218_not ; n2475
g2213 and n2474_not n2475_not ; n2476
g2214 and n2473 n2476 ; n2477
g2215 and n479 n2477_not ; n2478
g2216 and n2470_not n2478_not ; n2479
g2217 and n2462 n2479 ; n2480
g2218 and shift[6]_not n2480_not ; n2481
g2219 and n275 n1284_not ; n2482
g2220 and n288 n1301_not ; n2483
g2221 and n2482_not n2483_not ; n2484
g2222 and n302 n1349_not ; n2485
g2223 and n315 n1293_not ; n2486
g2224 and n2485_not n2486_not ; n2487
g2225 and n2484 n2487 ; n2488
g2226 and n479 n2488_not ; n2489
g2227 and n275 n1136_not ; n2490
g2228 and n288 n1153_not ; n2491
g2229 and n2490_not n2491_not ; n2492
g2230 and n302 n1276_not ; n2493
g2231 and n315 n1145_not ; n2494
g2232 and n2493_not n2494_not ; n2495
g2233 and n2492 n2495 ; n2496
g2234 and n426 n2496_not ; n2497
g2235 and n2489_not n2497_not ; n2498
g2236 and n275 n1357_not ; n2499
g2237 and n288 n1374_not ; n2500
g2238 and n2499_not n2500_not ; n2501
g2239 and n302 n1385_not ; n2502
g2240 and n315 n1366_not ; n2503
g2241 and n2502_not n2503_not ; n2504
g2242 and n2501 n2504 ; n2505
g2243 and n372 n2505_not ; n2506
g2244 and n275 n1393_not ; n2507
g2245 and n288 n1410_not ; n2508
g2246 and n2507_not n2508_not ; n2509
g2247 and n302 n1312_not ; n2510
g2248 and n315 n1402_not ; n2511
g2249 and n2510_not n2511_not ; n2512
g2250 and n2509 n2512 ; n2513
g2251 and n319 n2513_not ; n2514
g2252 and n2506_not n2514_not ; n2515
g2253 and n2498 n2515 ; n2516
g2254 and shift[6] n2516_not ; n2517
g2255 and n2481_not n2517_not ; result[14]
g2256 and n275 n1469_not ; n2519
g2257 and n288 n1486_not ; n2520
g2258 and n2519_not n2520_not ; n2521
g2259 and n302 n1534_not ; n2522
g2260 and n315 n1478_not ; n2523
g2261 and n2522_not n2523_not ; n2524
g2262 and n2521 n2524 ; n2525
g2263 and n319 n2525_not ; n2526
g2264 and n275 n1433_not ; n2527
g2265 and n288 n1450_not ; n2528
g2266 and n2527_not n2528_not ; n2529
g2267 and n302 n1461_not ; n2530
g2268 and n315 n1442_not ; n2531
g2269 and n2530_not n2531_not ; n2532
g2270 and n2529 n2532 ; n2533
g2271 and n372 n2533_not ; n2534
g2272 and n2526_not n2534_not ; n2535
g2273 and n275 n1654_not ; n2536
g2274 and n288 n1671_not ; n2537
g2275 and n2536_not n2537_not ; n2538
g2276 and n302 n1498_not ; n2539
g2277 and n315 n1663_not ; n2540
g2278 and n2539_not n2540_not ; n2541
g2279 and n2538 n2541 ; n2542
g2280 and n426 n2542_not ; n2543
g2281 and n275 n1506_not ; n2544
g2282 and n288 n1523_not ; n2545
g2283 and n2544_not n2545_not ; n2546
g2284 and n302 n1425_not ; n2547
g2285 and n315 n1515_not ; n2548
g2286 and n2547_not n2548_not ; n2549
g2287 and n2546 n2549 ; n2550
g2288 and n479 n2550_not ; n2551
g2289 and n2543_not n2551_not ; n2552
g2290 and n2535 n2552 ; n2553
g2291 and shift[6]_not n2553_not ; n2554
g2292 and n275 n1581_not ; n2555
g2293 and n288 n1598_not ; n2556
g2294 and n2555_not n2556_not ; n2557
g2295 and n302 n1609_not ; n2558
g2296 and n315 n1590_not ; n2559
g2297 and n2558_not n2559_not ; n2560
g2298 and n2557 n2560 ; n2561
g2299 and n479 n2561_not ; n2562
g2300 and n275 n1542_not ; n2563
g2301 and n288 n1559_not ; n2564
g2302 and n2563_not n2564_not ; n2565
g2303 and n302 n1573_not ; n2566
g2304 and n315 n1551_not ; n2567
g2305 and n2566_not n2567_not ; n2568
g2306 and n2565 n2568 ; n2569
g2307 and n426 n2569_not ; n2570
g2308 and n2562_not n2570_not ; n2571
g2309 and n275 n1617_not ; n2572
g2310 and n288 n1634_not ; n2573
g2311 and n2572_not n2573_not ; n2574
g2312 and n302 n1682_not ; n2575
g2313 and n315 n1626_not ; n2576
g2314 and n2575_not n2576_not ; n2577
g2315 and n2574 n2577 ; n2578
g2316 and n372 n2578_not ; n2579
g2317 and n275 n1690_not ; n2580
g2318 and n288 n1707_not ; n2581
g2319 and n2580_not n2581_not ; n2582
g2320 and n302 n1646_not ; n2583
g2321 and n315 n1699_not ; n2584
g2322 and n2583_not n2584_not ; n2585
g2323 and n2582 n2585 ; n2586
g2324 and n319 n2586_not ; n2587
g2325 and n2579_not n2587_not ; n2588
g2326 and n2571 n2588 ; n2589
g2327 and shift[6] n2589_not ; n2590
g2328 and n2554_not n2590_not ; result[15]
g2329 and n319 n371_not ; n2592
g2330 and n372 n478_not ; n2593
g2331 and n2592_not n2593_not ; n2594
g2332 and n426 n534_not ; n2595
g2333 and n425_not n479 ; n2596
g2334 and n2595_not n2596_not ; n2597
g2335 and n2594 n2597 ; n2598
g2336 and shift[6]_not n2598_not ; n2599
g2337 and n318_not n426 ; n2600
g2338 and n319 n586_not ; n2601
g2339 and n2600_not n2601_not ; n2602
g2340 and n479 n639_not ; n2603
g2341 and n372 n691_not ; n2604
g2342 and n2603_not n2604_not ; n2605
g2343 and n2602 n2605 ; n2606
g2344 and shift[6] n2606_not ; n2607
g2345 and n2599_not n2607_not ; result[16]
g2346 and n319 n799_not ; n2609
g2347 and n372 n904_not ; n2610
g2348 and n2609_not n2610_not ; n2611
g2349 and n426 n1011_not ; n2612
g2350 and n479 n852_not ; n2613
g2351 and n2612_not n2613_not ; n2614
g2352 and n2611 n2614 ; n2615
g2353 and shift[6]_not n2615_not ; n2616
g2354 and n479 n959_not ; n2617
g2355 and n426 n747_not ; n2618
g2356 and n2617_not n2618_not ; n2619
g2357 and n372 n1064_not ; n2620
g2358 and n319 n1116_not ; n2621
g2359 and n2620_not n2621_not ; n2622
g2360 and n2619 n2622 ; n2623
g2361 and shift[6] n2623_not ; n2624
g2362 and n2616_not n2624_not ; result[17]
g2363 and n319 n1192_not ; n2626
g2364 and n372 n1265_not ; n2627
g2365 and n2626_not n2627_not ; n2628
g2366 and n426 n1340_not ; n2629
g2367 and n479 n1229_not ; n2630
g2368 and n2629_not n2630_not ; n2631
g2369 and n2628 n2631 ; n2632
g2370 and shift[6]_not n2632_not ; n2633
g2371 and n479 n1304_not ; n2634
g2372 and n426 n1156_not ; n2635
g2373 and n2634_not n2635_not ; n2636
g2374 and n372 n1377_not ; n2637
g2375 and n319 n1413_not ; n2638
g2376 and n2637_not n2638_not ; n2639
g2377 and n2636 n2639 ; n2640
g2378 and shift[6] n2640_not ; n2641
g2379 and n2633_not n2641_not ; result[18]
g2380 and n372 n1453_not ; n2643
g2381 and n319 n1489_not ; n2644
g2382 and n2643_not n2644_not ; n2645
g2383 and n479 n1526_not ; n2646
g2384 and n426 n1674_not ; n2647
g2385 and n2646_not n2647_not ; n2648
g2386 and n2645 n2648 ; n2649
g2387 and shift[6]_not n2649_not ; n2650
g2388 and n479 n1601_not ; n2651
g2389 and n426 n1562_not ; n2652
g2390 and n2651_not n2652_not ; n2653
g2391 and n319 n1710_not ; n2654
g2392 and n372 n1637_not ; n2655
g2393 and n2654_not n2655_not ; n2656
g2394 and n2653 n2656 ; n2657
g2395 and shift[6] n2657_not ; n2658
g2396 and n2650_not n2658_not ; result[19]
g2397 and n319 n1730_not ; n2660
g2398 and n372 n1747_not ; n2661
g2399 and n2660_not n2661_not ; n2662
g2400 and n426 n1783_not ; n2663
g2401 and n479 n1739_not ; n2664
g2402 and n2663_not n2664_not ; n2665
g2403 and n2662 n2665 ; n2666
g2404 and shift[6]_not n2666_not ; n2667
g2405 and n426 n1722_not ; n2668
g2406 and n372 n1758_not ; n2669
g2407 and n2668_not n2669_not ; n2670
g2408 and n319 n1775_not ; n2671
g2409 and n479 n1766_not ; n2672
g2410 and n2671_not n2672_not ; n2673
g2411 and n2670 n2673 ; n2674
g2412 and shift[6] n2674_not ; n2675
g2413 and n2667_not n2675_not ; result[20]
g2414 and n319 n1803_not ; n2677
g2415 and n372 n1820_not ; n2678
g2416 and n2677_not n2678_not ; n2679
g2417 and n426 n1856_not ; n2680
g2418 and n479 n1812_not ; n2681
g2419 and n2680_not n2681_not ; n2682
g2420 and n2679 n2682 ; n2683
g2421 and shift[6]_not n2683_not ; n2684
g2422 and n426 n1795_not ; n2685
g2423 and n372 n1831_not ; n2686
g2424 and n2685_not n2686_not ; n2687
g2425 and n319 n1848_not ; n2688
g2426 and n479 n1839_not ; n2689
g2427 and n2688_not n2689_not ; n2690
g2428 and n2687 n2690 ; n2691
g2429 and shift[6] n2691_not ; n2692
g2430 and n2684_not n2692_not ; result[21]
g2431 and n319 n1876_not ; n2694
g2432 and n372 n1893_not ; n2695
g2433 and n2694_not n2695_not ; n2696
g2434 and n426 n1929_not ; n2697
g2435 and n479 n1885_not ; n2698
g2436 and n2697_not n2698_not ; n2699
g2437 and n2696 n2699 ; n2700
g2438 and shift[6]_not n2700_not ; n2701
g2439 and n426 n1868_not ; n2702
g2440 and n372 n1904_not ; n2703
g2441 and n2702_not n2703_not ; n2704
g2442 and n319 n1921_not ; n2705
g2443 and n479 n1912_not ; n2706
g2444 and n2705_not n2706_not ; n2707
g2445 and n2704 n2707 ; n2708
g2446 and shift[6] n2708_not ; n2709
g2447 and n2701_not n2709_not ; result[22]
g2448 and n319 n1949_not ; n2711
g2449 and n426 n2002_not ; n2712
g2450 and n2711_not n2712_not ; n2713
g2451 and n479 n1958_not ; n2714
g2452 and n372 n1966_not ; n2715
g2453 and n2714_not n2715_not ; n2716
g2454 and n2713 n2716 ; n2717
g2455 and shift[6]_not n2717_not ; n2718
g2456 and n372 n1977_not ; n2719
g2457 and n479 n1985_not ; n2720
g2458 and n2719_not n2720_not ; n2721
g2459 and n319 n1994_not ; n2722
g2460 and n426 n1941_not ; n2723
g2461 and n2722_not n2723_not ; n2724
g2462 and n2721 n2724 ; n2725
g2463 and shift[6] n2725_not ; n2726
g2464 and n2718_not n2726_not ; result[23]
g2465 and n319 n2022_not ; n2728
g2466 and n426 n2075_not ; n2729
g2467 and n2728_not n2729_not ; n2730
g2468 and n479 n2031_not ; n2731
g2469 and n372 n2039_not ; n2732
g2470 and n2731_not n2732_not ; n2733
g2471 and n2730 n2733 ; n2734
g2472 and shift[6]_not n2734_not ; n2735
g2473 and n372 n2050_not ; n2736
g2474 and n479 n2058_not ; n2737
g2475 and n2736_not n2737_not ; n2738
g2476 and n319 n2067_not ; n2739
g2477 and n426 n2014_not ; n2740
g2478 and n2739_not n2740_not ; n2741
g2479 and n2738 n2741 ; n2742
g2480 and shift[6] n2742_not ; n2743
g2481 and n2735_not n2743_not ; result[24]
g2482 and n319 n2095_not ; n2745
g2483 and n426 n2148_not ; n2746
g2484 and n2745_not n2746_not ; n2747
g2485 and n479 n2104_not ; n2748
g2486 and n372 n2112_not ; n2749
g2487 and n2748_not n2749_not ; n2750
g2488 and n2747 n2750 ; n2751
g2489 and shift[6]_not n2751_not ; n2752
g2490 and n372 n2123_not ; n2753
g2491 and n479 n2131_not ; n2754
g2492 and n2753_not n2754_not ; n2755
g2493 and n319 n2140_not ; n2756
g2494 and n426 n2087_not ; n2757
g2495 and n2756_not n2757_not ; n2758
g2496 and n2755 n2758 ; n2759
g2497 and shift[6] n2759_not ; n2760
g2498 and n2752_not n2760_not ; result[25]
g2499 and n319 n2168_not ; n2762
g2500 and n372 n2185_not ; n2763
g2501 and n2762_not n2763_not ; n2764
g2502 and n426 n2221_not ; n2765
g2503 and n479 n2177_not ; n2766
g2504 and n2765_not n2766_not ; n2767
g2505 and n2764 n2767 ; n2768
g2506 and shift[6]_not n2768_not ; n2769
g2507 and n372 n2196_not ; n2770
g2508 and n479 n2204_not ; n2771
g2509 and n2770_not n2771_not ; n2772
g2510 and n319 n2213_not ; n2773
g2511 and n426 n2160_not ; n2774
g2512 and n2773_not n2774_not ; n2775
g2513 and n2772 n2775 ; n2776
g2514 and shift[6] n2776_not ; n2777
g2515 and n2769_not n2777_not ; result[26]
g2516 and n319 n2241_not ; n2779
g2517 and n372 n2258_not ; n2780
g2518 and n2779_not n2780_not ; n2781
g2519 and n426 n2294_not ; n2782
g2520 and n479 n2250_not ; n2783
g2521 and n2782_not n2783_not ; n2784
g2522 and n2781 n2784 ; n2785
g2523 and shift[6]_not n2785_not ; n2786
g2524 and n372 n2269_not ; n2787
g2525 and n479 n2277_not ; n2788
g2526 and n2787_not n2788_not ; n2789
g2527 and n319 n2286_not ; n2790
g2528 and n426 n2233_not ; n2791
g2529 and n2790_not n2791_not ; n2792
g2530 and n2789 n2792 ; n2793
g2531 and shift[6] n2793_not ; n2794
g2532 and n2786_not n2794_not ; result[27]
g2533 and n319 n2314_not ; n2796
g2534 and n372 n2331_not ; n2797
g2535 and n2796_not n2797_not ; n2798
g2536 and n426 n2367_not ; n2799
g2537 and n479 n2323_not ; n2800
g2538 and n2799_not n2800_not ; n2801
g2539 and n2798 n2801 ; n2802
g2540 and shift[6]_not n2802_not ; n2803
g2541 and n372 n2342_not ; n2804
g2542 and n479 n2350_not ; n2805
g2543 and n2804_not n2805_not ; n2806
g2544 and n319 n2359_not ; n2807
g2545 and n426 n2306_not ; n2808
g2546 and n2807_not n2808_not ; n2809
g2547 and n2806 n2809 ; n2810
g2548 and shift[6] n2810_not ; n2811
g2549 and n2803_not n2811_not ; result[28]
g2550 and n319 n2387_not ; n2813
g2551 and n372 n2404_not ; n2814
g2552 and n2813_not n2814_not ; n2815
g2553 and n426 n2440_not ; n2816
g2554 and n479 n2396_not ; n2817
g2555 and n2816_not n2817_not ; n2818
g2556 and n2815 n2818 ; n2819
g2557 and shift[6]_not n2819_not ; n2820
g2558 and n372 n2415_not ; n2821
g2559 and n479 n2423_not ; n2822
g2560 and n2821_not n2822_not ; n2823
g2561 and n319 n2432_not ; n2824
g2562 and n426 n2379_not ; n2825
g2563 and n2824_not n2825_not ; n2826
g2564 and n2823 n2826 ; n2827
g2565 and shift[6] n2827_not ; n2828
g2566 and n2820_not n2828_not ; result[29]
g2567 and n319 n2460_not ; n2830
g2568 and n372 n2477_not ; n2831
g2569 and n2830_not n2831_not ; n2832
g2570 and n426 n2513_not ; n2833
g2571 and n479 n2469_not ; n2834
g2572 and n2833_not n2834_not ; n2835
g2573 and n2832 n2835 ; n2836
g2574 and shift[6]_not n2836_not ; n2837
g2575 and n372 n2488_not ; n2838
g2576 and n479 n2496_not ; n2839
g2577 and n2838_not n2839_not ; n2840
g2578 and n319 n2505_not ; n2841
g2579 and n426 n2452_not ; n2842
g2580 and n2841_not n2842_not ; n2843
g2581 and n2840 n2843 ; n2844
g2582 and shift[6] n2844_not ; n2845
g2583 and n2837_not n2845_not ; result[30]
g2584 and n319 n2533_not ; n2847
g2585 and n372 n2550_not ; n2848
g2586 and n2847_not n2848_not ; n2849
g2587 and n426 n2586_not ; n2850
g2588 and n479 n2542_not ; n2851
g2589 and n2850_not n2851_not ; n2852
g2590 and n2849 n2852 ; n2853
g2591 and shift[6]_not n2853_not ; n2854
g2592 and n372 n2561_not ; n2855
g2593 and n479 n2569_not ; n2856
g2594 and n2855_not n2856_not ; n2857
g2595 and n319 n2578_not ; n2858
g2596 and n426 n2525_not ; n2859
g2597 and n2858_not n2859_not ; n2860
g2598 and n2857 n2860 ; n2861
g2599 and shift[6] n2861_not ; n2862
g2600 and n2854_not n2862_not ; result[31]
g2601 and n319 n478_not ; n2864
g2602 and n372 n425_not ; n2865
g2603 and n2864_not n2865_not ; n2866
g2604 and n426 n586_not ; n2867
g2605 and n479 n534_not ; n2868
g2606 and n2867_not n2868_not ; n2869
g2607 and n2866 n2869 ; n2870
g2608 and shift[6]_not n2870_not ; n2871
g2609 and n318_not n479 ; n2872
g2610 and n371_not n426 ; n2873
g2611 and n2872_not n2873_not ; n2874
g2612 and n372 n639_not ; n2875
g2613 and n319 n691_not ; n2876
g2614 and n2875_not n2876_not ; n2877
g2615 and n2874 n2877 ; n2878
g2616 and shift[6] n2878_not ; n2879
g2617 and n2871_not n2879_not ; result[32]
g2618 and n319 n904_not ; n2881
g2619 and n372 n852_not ; n2882
g2620 and n2881_not n2882_not ; n2883
g2621 and n426 n1116_not ; n2884
g2622 and n479 n1011_not ; n2885
g2623 and n2884_not n2885_not ; n2886
g2624 and n2883 n2886 ; n2887
g2625 and shift[6]_not n2887_not ; n2888
g2626 and n372 n959_not ; n2889
g2627 and n479 n747_not ; n2890
g2628 and n2889_not n2890_not ; n2891
g2629 and n319 n1064_not ; n2892
g2630 and n426 n799_not ; n2893
g2631 and n2892_not n2893_not ; n2894
g2632 and n2891 n2894 ; n2895
g2633 and shift[6] n2895_not ; n2896
g2634 and n2888_not n2896_not ; result[33]
g2635 and n319 n1265_not ; n2898
g2636 and n372 n1229_not ; n2899
g2637 and n2898_not n2899_not ; n2900
g2638 and n426 n1413_not ; n2901
g2639 and n479 n1340_not ; n2902
g2640 and n2901_not n2902_not ; n2903
g2641 and n2900 n2903 ; n2904
g2642 and shift[6]_not n2904_not ; n2905
g2643 and n372 n1304_not ; n2906
g2644 and n479 n1156_not ; n2907
g2645 and n2906_not n2907_not ; n2908
g2646 and n319 n1377_not ; n2909
g2647 and n426 n1192_not ; n2910
g2648 and n2909_not n2910_not ; n2911
g2649 and n2908 n2911 ; n2912
g2650 and shift[6] n2912_not ; n2913
g2651 and n2905_not n2913_not ; result[34]
g2652 and n319 n1453_not ; n2915
g2653 and n426 n1710_not ; n2916
g2654 and n2915_not n2916_not ; n2917
g2655 and n372 n1526_not ; n2918
g2656 and n479 n1674_not ; n2919
g2657 and n2918_not n2919_not ; n2920
g2658 and n2917 n2920 ; n2921
g2659 and shift[6]_not n2921_not ; n2922
g2660 and n372 n1601_not ; n2923
g2661 and n426 n1489_not ; n2924
g2662 and n2923_not n2924_not ; n2925
g2663 and n319 n1637_not ; n2926
g2664 and n479 n1562_not ; n2927
g2665 and n2926_not n2927_not ; n2928
g2666 and n2925 n2928 ; n2929
g2667 and shift[6] n2929_not ; n2930
g2668 and n2922_not n2930_not ; result[35]
g2669 and n319 n1747_not ; n2932
g2670 and n372 n1739_not ; n2933
g2671 and n2932_not n2933_not ; n2934
g2672 and n426 n1775_not ; n2935
g2673 and n479 n1783_not ; n2936
g2674 and n2935_not n2936_not ; n2937
g2675 and n2934 n2937 ; n2938
g2676 and shift[6]_not n2938_not ; n2939
g2677 and n479 n1722_not ; n2940
g2678 and n426 n1730_not ; n2941
g2679 and n2940_not n2941_not ; n2942
g2680 and n372 n1766_not ; n2943
g2681 and n319 n1758_not ; n2944
g2682 and n2943_not n2944_not ; n2945
g2683 and n2942 n2945 ; n2946
g2684 and shift[6] n2946_not ; n2947
g2685 and n2939_not n2947_not ; result[36]
g2686 and n319 n1820_not ; n2949
g2687 and n372 n1812_not ; n2950
g2688 and n2949_not n2950_not ; n2951
g2689 and n426 n1848_not ; n2952
g2690 and n479 n1856_not ; n2953
g2691 and n2952_not n2953_not ; n2954
g2692 and n2951 n2954 ; n2955
g2693 and shift[6]_not n2955_not ; n2956
g2694 and n479 n1795_not ; n2957
g2695 and n426 n1803_not ; n2958
g2696 and n2957_not n2958_not ; n2959
g2697 and n372 n1839_not ; n2960
g2698 and n319 n1831_not ; n2961
g2699 and n2960_not n2961_not ; n2962
g2700 and n2959 n2962 ; n2963
g2701 and shift[6] n2963_not ; n2964
g2702 and n2956_not n2964_not ; result[37]
g2703 and n319 n1893_not ; n2966
g2704 and n372 n1885_not ; n2967
g2705 and n2966_not n2967_not ; n2968
g2706 and n426 n1921_not ; n2969
g2707 and n479 n1929_not ; n2970
g2708 and n2969_not n2970_not ; n2971
g2709 and n2968 n2971 ; n2972
g2710 and shift[6]_not n2972_not ; n2973
g2711 and n479 n1868_not ; n2974
g2712 and n426 n1876_not ; n2975
g2713 and n2974_not n2975_not ; n2976
g2714 and n372 n1912_not ; n2977
g2715 and n319 n1904_not ; n2978
g2716 and n2977_not n2978_not ; n2979
g2717 and n2976 n2979 ; n2980
g2718 and shift[6] n2980_not ; n2981
g2719 and n2973_not n2981_not ; result[38]
g2720 and n479 n2002_not ; n2983
g2721 and n426 n1994_not ; n2984
g2722 and n2983_not n2984_not ; n2985
g2723 and n372 n1958_not ; n2986
g2724 and n319 n1966_not ; n2987
g2725 and n2986_not n2987_not ; n2988
g2726 and n2985 n2988 ; n2989
g2727 and shift[6]_not n2989_not ; n2990
g2728 and n319 n1977_not ; n2991
g2729 and n372 n1985_not ; n2992
g2730 and n2991_not n2992_not ; n2993
g2731 and n426 n1949_not ; n2994
g2732 and n479 n1941_not ; n2995
g2733 and n2994_not n2995_not ; n2996
g2734 and n2993 n2996 ; n2997
g2735 and shift[6] n2997_not ; n2998
g2736 and n2990_not n2998_not ; result[39]
g2737 and n479 n2075_not ; n3000
g2738 and n426 n2067_not ; n3001
g2739 and n3000_not n3001_not ; n3002
g2740 and n372 n2031_not ; n3003
g2741 and n319 n2039_not ; n3004
g2742 and n3003_not n3004_not ; n3005
g2743 and n3002 n3005 ; n3006
g2744 and shift[6]_not n3006_not ; n3007
g2745 and n319 n2050_not ; n3008
g2746 and n372 n2058_not ; n3009
g2747 and n3008_not n3009_not ; n3010
g2748 and n426 n2022_not ; n3011
g2749 and n479 n2014_not ; n3012
g2750 and n3011_not n3012_not ; n3013
g2751 and n3010 n3013 ; n3014
g2752 and shift[6] n3014_not ; n3015
g2753 and n3007_not n3015_not ; result[40]
g2754 and n479 n2148_not ; n3017
g2755 and n426 n2140_not ; n3018
g2756 and n3017_not n3018_not ; n3019
g2757 and n372 n2104_not ; n3020
g2758 and n319 n2112_not ; n3021
g2759 and n3020_not n3021_not ; n3022
g2760 and n3019 n3022 ; n3023
g2761 and shift[6]_not n3023_not ; n3024
g2762 and n319 n2123_not ; n3025
g2763 and n372 n2131_not ; n3026
g2764 and n3025_not n3026_not ; n3027
g2765 and n426 n2095_not ; n3028
g2766 and n479 n2087_not ; n3029
g2767 and n3028_not n3029_not ; n3030
g2768 and n3027 n3030 ; n3031
g2769 and shift[6] n3031_not ; n3032
g2770 and n3024_not n3032_not ; result[41]
g2771 and n319 n2185_not ; n3034
g2772 and n372 n2177_not ; n3035
g2773 and n3034_not n3035_not ; n3036
g2774 and n426 n2213_not ; n3037
g2775 and n479 n2221_not ; n3038
g2776 and n3037_not n3038_not ; n3039
g2777 and n3036 n3039 ; n3040
g2778 and shift[6]_not n3040_not ; n3041
g2779 and n319 n2196_not ; n3042
g2780 and n372 n2204_not ; n3043
g2781 and n3042_not n3043_not ; n3044
g2782 and n426 n2168_not ; n3045
g2783 and n479 n2160_not ; n3046
g2784 and n3045_not n3046_not ; n3047
g2785 and n3044 n3047 ; n3048
g2786 and shift[6] n3048_not ; n3049
g2787 and n3041_not n3049_not ; result[42]
g2788 and n319 n2258_not ; n3051
g2789 and n372 n2250_not ; n3052
g2790 and n3051_not n3052_not ; n3053
g2791 and n426 n2286_not ; n3054
g2792 and n479 n2294_not ; n3055
g2793 and n3054_not n3055_not ; n3056
g2794 and n3053 n3056 ; n3057
g2795 and shift[6]_not n3057_not ; n3058
g2796 and n319 n2269_not ; n3059
g2797 and n372 n2277_not ; n3060
g2798 and n3059_not n3060_not ; n3061
g2799 and n426 n2241_not ; n3062
g2800 and n479 n2233_not ; n3063
g2801 and n3062_not n3063_not ; n3064
g2802 and n3061 n3064 ; n3065
g2803 and shift[6] n3065_not ; n3066
g2804 and n3058_not n3066_not ; result[43]
g2805 and n319 n2331_not ; n3068
g2806 and n372 n2323_not ; n3069
g2807 and n3068_not n3069_not ; n3070
g2808 and n426 n2359_not ; n3071
g2809 and n479 n2367_not ; n3072
g2810 and n3071_not n3072_not ; n3073
g2811 and n3070 n3073 ; n3074
g2812 and shift[6]_not n3074_not ; n3075
g2813 and n319 n2342_not ; n3076
g2814 and n372 n2350_not ; n3077
g2815 and n3076_not n3077_not ; n3078
g2816 and n426 n2314_not ; n3079
g2817 and n479 n2306_not ; n3080
g2818 and n3079_not n3080_not ; n3081
g2819 and n3078 n3081 ; n3082
g2820 and shift[6] n3082_not ; n3083
g2821 and n3075_not n3083_not ; result[44]
g2822 and n319 n2404_not ; n3085
g2823 and n372 n2396_not ; n3086
g2824 and n3085_not n3086_not ; n3087
g2825 and n426 n2432_not ; n3088
g2826 and n479 n2440_not ; n3089
g2827 and n3088_not n3089_not ; n3090
g2828 and n3087 n3090 ; n3091
g2829 and shift[6]_not n3091_not ; n3092
g2830 and n319 n2415_not ; n3093
g2831 and n372 n2423_not ; n3094
g2832 and n3093_not n3094_not ; n3095
g2833 and n426 n2387_not ; n3096
g2834 and n479 n2379_not ; n3097
g2835 and n3096_not n3097_not ; n3098
g2836 and n3095 n3098 ; n3099
g2837 and shift[6] n3099_not ; n3100
g2838 and n3092_not n3100_not ; result[45]
g2839 and n319 n2477_not ; n3102
g2840 and n372 n2469_not ; n3103
g2841 and n3102_not n3103_not ; n3104
g2842 and n426 n2505_not ; n3105
g2843 and n479 n2513_not ; n3106
g2844 and n3105_not n3106_not ; n3107
g2845 and n3104 n3107 ; n3108
g2846 and shift[6]_not n3108_not ; n3109
g2847 and n319 n2488_not ; n3110
g2848 and n372 n2496_not ; n3111
g2849 and n3110_not n3111_not ; n3112
g2850 and n426 n2460_not ; n3113
g2851 and n479 n2452_not ; n3114
g2852 and n3113_not n3114_not ; n3115
g2853 and n3112 n3115 ; n3116
g2854 and shift[6] n3116_not ; n3117
g2855 and n3109_not n3117_not ; result[46]
g2856 and n319 n2550_not ; n3119
g2857 and n372 n2542_not ; n3120
g2858 and n3119_not n3120_not ; n3121
g2859 and n426 n2578_not ; n3122
g2860 and n479 n2586_not ; n3123
g2861 and n3122_not n3123_not ; n3124
g2862 and n3121 n3124 ; n3125
g2863 and shift[6]_not n3125_not ; n3126
g2864 and n319 n2561_not ; n3127
g2865 and n372 n2569_not ; n3128
g2866 and n3127_not n3128_not ; n3129
g2867 and n426 n2533_not ; n3130
g2868 and n479 n2525_not ; n3131
g2869 and n3130_not n3131_not ; n3132
g2870 and n3129 n3132 ; n3133
g2871 and shift[6] n3133_not ; n3134
g2872 and n3126_not n3134_not ; result[47]
g2873 and n319 n425_not ; n3136
g2874 and n372 n534_not ; n3137
g2875 and n3136_not n3137_not ; n3138
g2876 and n426 n691_not ; n3139
g2877 and n479 n586_not ; n3140
g2878 and n3139_not n3140_not ; n3141
g2879 and n3138 n3141 ; n3142
g2880 and shift[6]_not n3142_not ; n3143
g2881 and n318_not n372 ; n3144
g2882 and n371_not n479 ; n3145
g2883 and n3144_not n3145_not ; n3146
g2884 and n319 n639_not ; n3147
g2885 and n426 n478_not ; n3148
g2886 and n3147_not n3148_not ; n3149
g2887 and n3146 n3149 ; n3150
g2888 and shift[6] n3150_not ; n3151
g2889 and n3143_not n3151_not ; result[48]
g2890 and n319 n852_not ; n3153
g2891 and n372 n1011_not ; n3154
g2892 and n3153_not n3154_not ; n3155
g2893 and n426 n1064_not ; n3156
g2894 and n479 n1116_not ; n3157
g2895 and n3156_not n3157_not ; n3158
g2896 and n3155 n3158 ; n3159
g2897 and shift[6]_not n3159_not ; n3160
g2898 and n319 n959_not ; n3161
g2899 and n372 n747_not ; n3162
g2900 and n3161_not n3162_not ; n3163
g2901 and n426 n904_not ; n3164
g2902 and n479 n799_not ; n3165
g2903 and n3164_not n3165_not ; n3166
g2904 and n3163 n3166 ; n3167
g2905 and shift[6] n3167_not ; n3168
g2906 and n3160_not n3168_not ; result[49]
g2907 and n319 n1229_not ; n3170
g2908 and n372 n1340_not ; n3171
g2909 and n3170_not n3171_not ; n3172
g2910 and n426 n1377_not ; n3173
g2911 and n479 n1413_not ; n3174
g2912 and n3173_not n3174_not ; n3175
g2913 and n3172 n3175 ; n3176
g2914 and shift[6]_not n3176_not ; n3177
g2915 and n319 n1304_not ; n3178
g2916 and n372 n1156_not ; n3179
g2917 and n3178_not n3179_not ; n3180
g2918 and n426 n1265_not ; n3181
g2919 and n479 n1192_not ; n3182
g2920 and n3181_not n3182_not ; n3183
g2921 and n3180 n3183 ; n3184
g2922 and shift[6] n3184_not ; n3185
g2923 and n3177_not n3185_not ; result[50]
g2924 and n426 n1637_not ; n3187
g2925 and n479 n1710_not ; n3188
g2926 and n3187_not n3188_not ; n3189
g2927 and n319 n1526_not ; n3190
g2928 and n372 n1674_not ; n3191
g2929 and n3190_not n3191_not ; n3192
g2930 and n3189 n3192 ; n3193
g2931 and shift[6]_not n3193_not ; n3194
g2932 and n319 n1601_not ; n3195
g2933 and n426 n1453_not ; n3196
g2934 and n3195_not n3196_not ; n3197
g2935 and n372 n1562_not ; n3198
g2936 and n479 n1489_not ; n3199
g2937 and n3198_not n3199_not ; n3200
g2938 and n3197 n3200 ; n3201
g2939 and shift[6] n3201_not ; n3202
g2940 and n3194_not n3202_not ; result[51]
g2941 and n426 n1758_not ; n3204
g2942 and n319 n1739_not ; n3205
g2943 and n3204_not n3205_not ; n3206
g2944 and n479 n1775_not ; n3207
g2945 and n372 n1783_not ; n3208
g2946 and n3207_not n3208_not ; n3209
g2947 and n3206 n3209 ; n3210
g2948 and shift[6]_not n3210_not ; n3211
g2949 and n372 n1722_not ; n3212
g2950 and n479 n1730_not ; n3213
g2951 and n3212_not n3213_not ; n3214
g2952 and n426 n1747_not ; n3215
g2953 and n319 n1766_not ; n3216
g2954 and n3215_not n3216_not ; n3217
g2955 and n3214 n3217 ; n3218
g2956 and shift[6] n3218_not ; n3219
g2957 and n3211_not n3219_not ; result[52]
g2958 and n426 n1831_not ; n3221
g2959 and n319 n1812_not ; n3222
g2960 and n3221_not n3222_not ; n3223
g2961 and n479 n1848_not ; n3224
g2962 and n372 n1856_not ; n3225
g2963 and n3224_not n3225_not ; n3226
g2964 and n3223 n3226 ; n3227
g2965 and shift[6]_not n3227_not ; n3228
g2966 and n372 n1795_not ; n3229
g2967 and n479 n1803_not ; n3230
g2968 and n3229_not n3230_not ; n3231
g2969 and n426 n1820_not ; n3232
g2970 and n319 n1839_not ; n3233
g2971 and n3232_not n3233_not ; n3234
g2972 and n3231 n3234 ; n3235
g2973 and shift[6] n3235_not ; n3236
g2974 and n3228_not n3236_not ; result[53]
g2975 and n426 n1904_not ; n3238
g2976 and n319 n1885_not ; n3239
g2977 and n3238_not n3239_not ; n3240
g2978 and n479 n1921_not ; n3241
g2979 and n372 n1929_not ; n3242
g2980 and n3241_not n3242_not ; n3243
g2981 and n3240 n3243 ; n3244
g2982 and shift[6]_not n3244_not ; n3245
g2983 and n372 n1868_not ; n3246
g2984 and n479 n1876_not ; n3247
g2985 and n3246_not n3247_not ; n3248
g2986 and n426 n1893_not ; n3249
g2987 and n319 n1912_not ; n3250
g2988 and n3249_not n3250_not ; n3251
g2989 and n3248 n3251 ; n3252
g2990 and shift[6] n3252_not ; n3253
g2991 and n3245_not n3253_not ; result[54]
g2992 and n426 n1977_not ; n3255
g2993 and n372 n2002_not ; n3256
g2994 and n3255_not n3256_not ; n3257
g2995 and n319 n1958_not ; n3258
g2996 and n479 n1994_not ; n3259
g2997 and n3258_not n3259_not ; n3260
g2998 and n3257 n3260 ; n3261
g2999 and shift[6]_not n3261_not ; n3262
g3000 and n319 n1985_not ; n3263
g3001 and n372 n1941_not ; n3264
g3002 and n3263_not n3264_not ; n3265
g3003 and n426 n1966_not ; n3266
g3004 and n479 n1949_not ; n3267
g3005 and n3266_not n3267_not ; n3268
g3006 and n3265 n3268 ; n3269
g3007 and shift[6] n3269_not ; n3270
g3008 and n3262_not n3270_not ; result[55]
g3009 and n426 n2050_not ; n3272
g3010 and n372 n2075_not ; n3273
g3011 and n3272_not n3273_not ; n3274
g3012 and n319 n2031_not ; n3275
g3013 and n479 n2067_not ; n3276
g3014 and n3275_not n3276_not ; n3277
g3015 and n3274 n3277 ; n3278
g3016 and shift[6]_not n3278_not ; n3279
g3017 and n319 n2058_not ; n3280
g3018 and n372 n2014_not ; n3281
g3019 and n3280_not n3281_not ; n3282
g3020 and n426 n2039_not ; n3283
g3021 and n479 n2022_not ; n3284
g3022 and n3283_not n3284_not ; n3285
g3023 and n3282 n3285 ; n3286
g3024 and shift[6] n3286_not ; n3287
g3025 and n3279_not n3287_not ; result[56]
g3026 and n426 n2123_not ; n3289
g3027 and n372 n2148_not ; n3290
g3028 and n3289_not n3290_not ; n3291
g3029 and n319 n2104_not ; n3292
g3030 and n479 n2140_not ; n3293
g3031 and n3292_not n3293_not ; n3294
g3032 and n3291 n3294 ; n3295
g3033 and shift[6]_not n3295_not ; n3296
g3034 and n319 n2131_not ; n3297
g3035 and n372 n2087_not ; n3298
g3036 and n3297_not n3298_not ; n3299
g3037 and n426 n2112_not ; n3300
g3038 and n479 n2095_not ; n3301
g3039 and n3300_not n3301_not ; n3302
g3040 and n3299 n3302 ; n3303
g3041 and shift[6] n3303_not ; n3304
g3042 and n3296_not n3304_not ; result[57]
g3043 and n426 n2196_not ; n3306
g3044 and n319 n2177_not ; n3307
g3045 and n3306_not n3307_not ; n3308
g3046 and n479 n2213_not ; n3309
g3047 and n372 n2221_not ; n3310
g3048 and n3309_not n3310_not ; n3311
g3049 and n3308 n3311 ; n3312
g3050 and shift[6]_not n3312_not ; n3313
g3051 and n319 n2204_not ; n3314
g3052 and n372 n2160_not ; n3315
g3053 and n3314_not n3315_not ; n3316
g3054 and n426 n2185_not ; n3317
g3055 and n479 n2168_not ; n3318
g3056 and n3317_not n3318_not ; n3319
g3057 and n3316 n3319 ; n3320
g3058 and shift[6] n3320_not ; n3321
g3059 and n3313_not n3321_not ; result[58]
g3060 and n426 n2269_not ; n3323
g3061 and n319 n2250_not ; n3324
g3062 and n3323_not n3324_not ; n3325
g3063 and n479 n2286_not ; n3326
g3064 and n372 n2294_not ; n3327
g3065 and n3326_not n3327_not ; n3328
g3066 and n3325 n3328 ; n3329
g3067 and shift[6]_not n3329_not ; n3330
g3068 and n319 n2277_not ; n3331
g3069 and n372 n2233_not ; n3332
g3070 and n3331_not n3332_not ; n3333
g3071 and n426 n2258_not ; n3334
g3072 and n479 n2241_not ; n3335
g3073 and n3334_not n3335_not ; n3336
g3074 and n3333 n3336 ; n3337
g3075 and shift[6] n3337_not ; n3338
g3076 and n3330_not n3338_not ; result[59]
g3077 and n426 n2342_not ; n3340
g3078 and n319 n2323_not ; n3341
g3079 and n3340_not n3341_not ; n3342
g3080 and n479 n2359_not ; n3343
g3081 and n372 n2367_not ; n3344
g3082 and n3343_not n3344_not ; n3345
g3083 and n3342 n3345 ; n3346
g3084 and shift[6]_not n3346_not ; n3347
g3085 and n319 n2350_not ; n3348
g3086 and n372 n2306_not ; n3349
g3087 and n3348_not n3349_not ; n3350
g3088 and n426 n2331_not ; n3351
g3089 and n479 n2314_not ; n3352
g3090 and n3351_not n3352_not ; n3353
g3091 and n3350 n3353 ; n3354
g3092 and shift[6] n3354_not ; n3355
g3093 and n3347_not n3355_not ; result[60]
g3094 and n426 n2415_not ; n3357
g3095 and n319 n2396_not ; n3358
g3096 and n3357_not n3358_not ; n3359
g3097 and n479 n2432_not ; n3360
g3098 and n372 n2440_not ; n3361
g3099 and n3360_not n3361_not ; n3362
g3100 and n3359 n3362 ; n3363
g3101 and shift[6]_not n3363_not ; n3364
g3102 and n319 n2423_not ; n3365
g3103 and n372 n2379_not ; n3366
g3104 and n3365_not n3366_not ; n3367
g3105 and n426 n2404_not ; n3368
g3106 and n479 n2387_not ; n3369
g3107 and n3368_not n3369_not ; n3370
g3108 and n3367 n3370 ; n3371
g3109 and shift[6] n3371_not ; n3372
g3110 and n3364_not n3372_not ; result[61]
g3111 and n426 n2488_not ; n3374
g3112 and n319 n2469_not ; n3375
g3113 and n3374_not n3375_not ; n3376
g3114 and n479 n2505_not ; n3377
g3115 and n372 n2513_not ; n3378
g3116 and n3377_not n3378_not ; n3379
g3117 and n3376 n3379 ; n3380
g3118 and shift[6]_not n3380_not ; n3381
g3119 and n319 n2496_not ; n3382
g3120 and n372 n2452_not ; n3383
g3121 and n3382_not n3383_not ; n3384
g3122 and n426 n2477_not ; n3385
g3123 and n479 n2460_not ; n3386
g3124 and n3385_not n3386_not ; n3387
g3125 and n3384 n3387 ; n3388
g3126 and shift[6] n3388_not ; n3389
g3127 and n3381_not n3389_not ; result[62]
g3128 and n426 n2561_not ; n3391
g3129 and n319 n2542_not ; n3392
g3130 and n3391_not n3392_not ; n3393
g3131 and n479 n2578_not ; n3394
g3132 and n372 n2586_not ; n3395
g3133 and n3394_not n3395_not ; n3396
g3134 and n3393 n3396 ; n3397
g3135 and shift[6]_not n3397_not ; n3398
g3136 and n319 n2569_not ; n3399
g3137 and n372 n2525_not ; n3400
g3138 and n3399_not n3400_not ; n3401
g3139 and n426 n2550_not ; n3402
g3140 and n479 n2533_not ; n3403
g3141 and n3402_not n3403_not ; n3404
g3142 and n3401 n3404 ; n3405
g3143 and shift[6] n3405_not ; n3406
g3144 and n3398_not n3406_not ; result[63]
g3145 and shift[6]_not n694_not ; n3408
g3146 and shift[6] n482_not ; n3409
g3147 and n3408_not n3409_not ; result[64]
g3148 and shift[6]_not n1119_not ; n3411
g3149 and shift[6] n907_not ; n3412
g3150 and n3411_not n3412_not ; result[65]
g3151 and shift[6]_not n1416_not ; n3414
g3152 and shift[6] n1268_not ; n3415
g3153 and n3414_not n3415_not ; result[66]
g3154 and shift[6]_not n1713_not ; n3417
g3155 and shift[6] n1565_not ; n3418
g3156 and n3417_not n3418_not ; result[67]
g3157 and shift[6]_not n1786_not ; n3420
g3158 and shift[6] n1750_not ; n3421
g3159 and n3420_not n3421_not ; result[68]
g3160 and shift[6]_not n1859_not ; n3423
g3161 and shift[6] n1823_not ; n3424
g3162 and n3423_not n3424_not ; result[69]
g3163 and shift[6]_not n1932_not ; n3426
g3164 and shift[6] n1896_not ; n3427
g3165 and n3426_not n3427_not ; result[70]
g3166 and shift[6]_not n2005_not ; n3429
g3167 and shift[6] n1969_not ; n3430
g3168 and n3429_not n3430_not ; result[71]
g3169 and shift[6]_not n2078_not ; n3432
g3170 and shift[6] n2042_not ; n3433
g3171 and n3432_not n3433_not ; result[72]
g3172 and shift[6]_not n2151_not ; n3435
g3173 and shift[6] n2115_not ; n3436
g3174 and n3435_not n3436_not ; result[73]
g3175 and shift[6]_not n2224_not ; n3438
g3176 and shift[6] n2188_not ; n3439
g3177 and n3438_not n3439_not ; result[74]
g3178 and shift[6]_not n2297_not ; n3441
g3179 and shift[6] n2261_not ; n3442
g3180 and n3441_not n3442_not ; result[75]
g3181 and shift[6]_not n2370_not ; n3444
g3182 and shift[6] n2334_not ; n3445
g3183 and n3444_not n3445_not ; result[76]
g3184 and shift[6]_not n2443_not ; n3447
g3185 and shift[6] n2407_not ; n3448
g3186 and n3447_not n3448_not ; result[77]
g3187 and shift[6]_not n2516_not ; n3450
g3188 and shift[6] n2480_not ; n3451
g3189 and n3450_not n3451_not ; result[78]
g3190 and shift[6]_not n2589_not ; n3453
g3191 and shift[6] n2553_not ; n3454
g3192 and n3453_not n3454_not ; result[79]
g3193 and shift[6]_not n2606_not ; n3456
g3194 and shift[6] n2598_not ; n3457
g3195 and n3456_not n3457_not ; result[80]
g3196 and shift[6]_not n2623_not ; n3459
g3197 and shift[6] n2615_not ; n3460
g3198 and n3459_not n3460_not ; result[81]
g3199 and shift[6]_not n2640_not ; n3462
g3200 and shift[6] n2632_not ; n3463
g3201 and n3462_not n3463_not ; result[82]
g3202 and shift[6]_not n2657_not ; n3465
g3203 and shift[6] n2649_not ; n3466
g3204 and n3465_not n3466_not ; result[83]
g3205 and shift[6]_not n2674_not ; n3468
g3206 and shift[6] n2666_not ; n3469
g3207 and n3468_not n3469_not ; result[84]
g3208 and shift[6]_not n2691_not ; n3471
g3209 and shift[6] n2683_not ; n3472
g3210 and n3471_not n3472_not ; result[85]
g3211 and shift[6]_not n2708_not ; n3474
g3212 and shift[6] n2700_not ; n3475
g3213 and n3474_not n3475_not ; result[86]
g3214 and shift[6]_not n2725_not ; n3477
g3215 and shift[6] n2717_not ; n3478
g3216 and n3477_not n3478_not ; result[87]
g3217 and shift[6]_not n2742_not ; n3480
g3218 and shift[6] n2734_not ; n3481
g3219 and n3480_not n3481_not ; result[88]
g3220 and shift[6]_not n2759_not ; n3483
g3221 and shift[6] n2751_not ; n3484
g3222 and n3483_not n3484_not ; result[89]
g3223 and shift[6]_not n2776_not ; n3486
g3224 and shift[6] n2768_not ; n3487
g3225 and n3486_not n3487_not ; result[90]
g3226 and shift[6]_not n2793_not ; n3489
g3227 and shift[6] n2785_not ; n3490
g3228 and n3489_not n3490_not ; result[91]
g3229 and shift[6]_not n2810_not ; n3492
g3230 and shift[6] n2802_not ; n3493
g3231 and n3492_not n3493_not ; result[92]
g3232 and shift[6]_not n2827_not ; n3495
g3233 and shift[6] n2819_not ; n3496
g3234 and n3495_not n3496_not ; result[93]
g3235 and shift[6]_not n2844_not ; n3498
g3236 and shift[6] n2836_not ; n3499
g3237 and n3498_not n3499_not ; result[94]
g3238 and shift[6]_not n2861_not ; n3501
g3239 and shift[6] n2853_not ; n3502
g3240 and n3501_not n3502_not ; result[95]
g3241 and shift[6]_not n2878_not ; n3504
g3242 and shift[6] n2870_not ; n3505
g3243 and n3504_not n3505_not ; result[96]
g3244 and shift[6]_not n2895_not ; n3507
g3245 and shift[6] n2887_not ; n3508
g3246 and n3507_not n3508_not ; result[97]
g3247 and shift[6]_not n2912_not ; n3510
g3248 and shift[6] n2904_not ; n3511
g3249 and n3510_not n3511_not ; result[98]
g3250 and shift[6]_not n2929_not ; n3513
g3251 and shift[6] n2921_not ; n3514
g3252 and n3513_not n3514_not ; result[99]
g3253 and shift[6]_not n2946_not ; n3516
g3254 and shift[6] n2938_not ; n3517
g3255 and n3516_not n3517_not ; result[100]
g3256 and shift[6]_not n2963_not ; n3519
g3257 and shift[6] n2955_not ; n3520
g3258 and n3519_not n3520_not ; result[101]
g3259 and shift[6]_not n2980_not ; n3522
g3260 and shift[6] n2972_not ; n3523
g3261 and n3522_not n3523_not ; result[102]
g3262 and shift[6]_not n2997_not ; n3525
g3263 and shift[6] n2989_not ; n3526
g3264 and n3525_not n3526_not ; result[103]
g3265 and shift[6]_not n3014_not ; n3528
g3266 and shift[6] n3006_not ; n3529
g3267 and n3528_not n3529_not ; result[104]
g3268 and shift[6]_not n3031_not ; n3531
g3269 and shift[6] n3023_not ; n3532
g3270 and n3531_not n3532_not ; result[105]
g3271 and shift[6]_not n3048_not ; n3534
g3272 and shift[6] n3040_not ; n3535
g3273 and n3534_not n3535_not ; result[106]
g3274 and shift[6]_not n3065_not ; n3537
g3275 and shift[6] n3057_not ; n3538
g3276 and n3537_not n3538_not ; result[107]
g3277 and shift[6]_not n3082_not ; n3540
g3278 and shift[6] n3074_not ; n3541
g3279 and n3540_not n3541_not ; result[108]
g3280 and shift[6]_not n3099_not ; n3543
g3281 and shift[6] n3091_not ; n3544
g3282 and n3543_not n3544_not ; result[109]
g3283 and shift[6]_not n3116_not ; n3546
g3284 and shift[6] n3108_not ; n3547
g3285 and n3546_not n3547_not ; result[110]
g3286 and shift[6]_not n3133_not ; n3549
g3287 and shift[6] n3125_not ; n3550
g3288 and n3549_not n3550_not ; result[111]
g3289 and shift[6]_not n3150_not ; n3552
g3290 and shift[6] n3142_not ; n3553
g3291 and n3552_not n3553_not ; result[112]
g3292 and shift[6]_not n3167_not ; n3555
g3293 and shift[6] n3159_not ; n3556
g3294 and n3555_not n3556_not ; result[113]
g3295 and shift[6]_not n3184_not ; n3558
g3296 and shift[6] n3176_not ; n3559
g3297 and n3558_not n3559_not ; result[114]
g3298 and shift[6]_not n3201_not ; n3561
g3299 and shift[6] n3193_not ; n3562
g3300 and n3561_not n3562_not ; result[115]
g3301 and shift[6]_not n3218_not ; n3564
g3302 and shift[6] n3210_not ; n3565
g3303 and n3564_not n3565_not ; result[116]
g3304 and shift[6]_not n3235_not ; n3567
g3305 and shift[6] n3227_not ; n3568
g3306 and n3567_not n3568_not ; result[117]
g3307 and shift[6]_not n3252_not ; n3570
g3308 and shift[6] n3244_not ; n3571
g3309 and n3570_not n3571_not ; result[118]
g3310 and shift[6]_not n3269_not ; n3573
g3311 and shift[6] n3261_not ; n3574
g3312 and n3573_not n3574_not ; result[119]
g3313 and shift[6]_not n3286_not ; n3576
g3314 and shift[6] n3278_not ; n3577
g3315 and n3576_not n3577_not ; result[120]
g3316 and shift[6]_not n3303_not ; n3579
g3317 and shift[6] n3295_not ; n3580
g3318 and n3579_not n3580_not ; result[121]
g3319 and shift[6]_not n3320_not ; n3582
g3320 and shift[6] n3312_not ; n3583
g3321 and n3582_not n3583_not ; result[122]
g3322 and shift[6]_not n3337_not ; n3585
g3323 and shift[6] n3329_not ; n3586
g3324 and n3585_not n3586_not ; result[123]
g3325 and shift[6]_not n3354_not ; n3588
g3326 and shift[6] n3346_not ; n3589
g3327 and n3588_not n3589_not ; result[124]
g3328 and shift[6]_not n3371_not ; n3591
g3329 and shift[6] n3363_not ; n3592
g3330 and n3591_not n3592_not ; result[125]
g3331 and shift[6]_not n3388_not ; n3594
g3332 and shift[6] n3380_not ; n3595
g3333 and n3594_not n3595_not ; result[126]
g3334 and shift[6]_not n3405_not ; n3597
g3335 and shift[6] n3397_not ; n3598
g3336 and n3597_not n3598_not ; result[127]
g3337 not shift[0] ; shift[0]_not
g3338 not n265 ; n265_not
g3339 not n267 ; n267_not
g3340 not shift[1] ; shift[1]_not
g3341 not n270 ; n270_not
g3342 not n272 ; n272_not
g3343 not shift[2] ; shift[2]_not
g3344 not shift[3] ; shift[3]_not
g3345 not n274 ; n274_not
g3346 not n278 ; n278_not
g3347 not n280 ; n280_not
g3348 not n283 ; n283_not
g3349 not n285 ; n285_not
g3350 not n287 ; n287_not
g3351 not n276 ; n276_not
g3352 not n289 ; n289_not
g3353 not n292 ; n292_not
g3354 not n294 ; n294_not
g3355 not n297 ; n297_not
g3356 not n299 ; n299_not
g3357 not n301 ; n301_not
g3358 not n305 ; n305_not
g3359 not n307 ; n307_not
g3360 not n310 ; n310_not
g3361 not n312 ; n312_not
g3362 not n314 ; n314_not
g3363 not n303 ; n303_not
g3364 not n316 ; n316_not
g3365 not n318 ; n318_not
g3366 not n322 ; n322_not
g3367 not n324 ; n324_not
g3368 not n327 ; n327_not
g3369 not n329 ; n329_not
g3370 not n331 ; n331_not
g3371 not n334 ; n334_not
g3372 not n336 ; n336_not
g3373 not n339 ; n339_not
g3374 not n341 ; n341_not
g3375 not n343 ; n343_not
g3376 not n332 ; n332_not
g3377 not n344 ; n344_not
g3378 not n347 ; n347_not
g3379 not n349 ; n349_not
g3380 not n352 ; n352_not
g3381 not n354 ; n354_not
g3382 not n356 ; n356_not
g3383 not n359 ; n359_not
g3384 not n361 ; n361_not
g3385 not n364 ; n364_not
g3386 not n366 ; n366_not
g3387 not n368 ; n368_not
g3388 not n357 ; n357_not
g3389 not n369 ; n369_not
g3390 not shift[4] ; shift[4]_not
g3391 not n371 ; n371_not
g3392 not n320 ; n320_not
g3393 not n373 ; n373_not
g3394 not n376 ; n376_not
g3395 not n378 ; n378_not
g3396 not n381 ; n381_not
g3397 not n383 ; n383_not
g3398 not n385 ; n385_not
g3399 not n388 ; n388_not
g3400 not n390 ; n390_not
g3401 not n393 ; n393_not
g3402 not n395 ; n395_not
g3403 not n397 ; n397_not
g3404 not n386 ; n386_not
g3405 not n398 ; n398_not
g3406 not n401 ; n401_not
g3407 not n403 ; n403_not
g3408 not n406 ; n406_not
g3409 not n408 ; n408_not
g3410 not n410 ; n410_not
g3411 not n413 ; n413_not
g3412 not n415 ; n415_not
g3413 not n418 ; n418_not
g3414 not n420 ; n420_not
g3415 not n422 ; n422_not
g3416 not n411 ; n411_not
g3417 not n423 ; n423_not
g3418 not shift[5] ; shift[5]_not
g3419 not n425 ; n425_not
g3420 not n429 ; n429_not
g3421 not n431 ; n431_not
g3422 not n434 ; n434_not
g3423 not n436 ; n436_not
g3424 not n438 ; n438_not
g3425 not n441 ; n441_not
g3426 not n443 ; n443_not
g3427 not n446 ; n446_not
g3428 not n448 ; n448_not
g3429 not n450 ; n450_not
g3430 not n439 ; n439_not
g3431 not n451 ; n451_not
g3432 not n454 ; n454_not
g3433 not n456 ; n456_not
g3434 not n459 ; n459_not
g3435 not n461 ; n461_not
g3436 not n463 ; n463_not
g3437 not n466 ; n466_not
g3438 not n468 ; n468_not
g3439 not n471 ; n471_not
g3440 not n473 ; n473_not
g3441 not n475 ; n475_not
g3442 not n464 ; n464_not
g3443 not n476 ; n476_not
g3444 not n478 ; n478_not
g3445 not n427 ; n427_not
g3446 not n480 ; n480_not
g3447 not shift[6] ; shift[6]_not
g3448 not n482 ; n482_not
g3449 not n485 ; n485_not
g3450 not n487 ; n487_not
g3451 not n490 ; n490_not
g3452 not n492 ; n492_not
g3453 not n494 ; n494_not
g3454 not n497 ; n497_not
g3455 not n499 ; n499_not
g3456 not n502 ; n502_not
g3457 not n504 ; n504_not
g3458 not n506 ; n506_not
g3459 not n495 ; n495_not
g3460 not n507 ; n507_not
g3461 not n510 ; n510_not
g3462 not n512 ; n512_not
g3463 not n515 ; n515_not
g3464 not n517 ; n517_not
g3465 not n519 ; n519_not
g3466 not n522 ; n522_not
g3467 not n524 ; n524_not
g3468 not n527 ; n527_not
g3469 not n529 ; n529_not
g3470 not n531 ; n531_not
g3471 not n520 ; n520_not
g3472 not n532 ; n532_not
g3473 not n534 ; n534_not
g3474 not n537 ; n537_not
g3475 not n539 ; n539_not
g3476 not n542 ; n542_not
g3477 not n544 ; n544_not
g3478 not n546 ; n546_not
g3479 not n549 ; n549_not
g3480 not n551 ; n551_not
g3481 not n554 ; n554_not
g3482 not n556 ; n556_not
g3483 not n558 ; n558_not
g3484 not n547 ; n547_not
g3485 not n559 ; n559_not
g3486 not n562 ; n562_not
g3487 not n564 ; n564_not
g3488 not n567 ; n567_not
g3489 not n569 ; n569_not
g3490 not n571 ; n571_not
g3491 not n574 ; n574_not
g3492 not n576 ; n576_not
g3493 not n579 ; n579_not
g3494 not n581 ; n581_not
g3495 not n583 ; n583_not
g3496 not n572 ; n572_not
g3497 not n584 ; n584_not
g3498 not n586 ; n586_not
g3499 not n535 ; n535_not
g3500 not n587 ; n587_not
g3501 not n590 ; n590_not
g3502 not n592 ; n592_not
g3503 not n595 ; n595_not
g3504 not n597 ; n597_not
g3505 not n599 ; n599_not
g3506 not n602 ; n602_not
g3507 not n604 ; n604_not
g3508 not n607 ; n607_not
g3509 not n609 ; n609_not
g3510 not n611 ; n611_not
g3511 not n600 ; n600_not
g3512 not n612 ; n612_not
g3513 not n615 ; n615_not
g3514 not n617 ; n617_not
g3515 not n620 ; n620_not
g3516 not n622 ; n622_not
g3517 not n624 ; n624_not
g3518 not n627 ; n627_not
g3519 not n629 ; n629_not
g3520 not n632 ; n632_not
g3521 not n634 ; n634_not
g3522 not n636 ; n636_not
g3523 not n625 ; n625_not
g3524 not n637 ; n637_not
g3525 not n639 ; n639_not
g3526 not n642 ; n642_not
g3527 not n644 ; n644_not
g3528 not n647 ; n647_not
g3529 not n649 ; n649_not
g3530 not n651 ; n651_not
g3531 not n654 ; n654_not
g3532 not n656 ; n656_not
g3533 not n659 ; n659_not
g3534 not n661 ; n661_not
g3535 not n663 ; n663_not
g3536 not n652 ; n652_not
g3537 not n664 ; n664_not
g3538 not n667 ; n667_not
g3539 not n669 ; n669_not
g3540 not n672 ; n672_not
g3541 not n674 ; n674_not
g3542 not n676 ; n676_not
g3543 not n679 ; n679_not
g3544 not n681 ; n681_not
g3545 not n684 ; n684_not
g3546 not n686 ; n686_not
g3547 not n688 ; n688_not
g3548 not n677 ; n677_not
g3549 not n689 ; n689_not
g3550 not n691 ; n691_not
g3551 not n640 ; n640_not
g3552 not n692 ; n692_not
g3553 not n694 ; n694_not
g3554 not n483 ; n483_not
g3555 not n695 ; n695_not
g3556 not n698 ; n698_not
g3557 not n700 ; n700_not
g3558 not n703 ; n703_not
g3559 not n705 ; n705_not
g3560 not n707 ; n707_not
g3561 not n710 ; n710_not
g3562 not n712 ; n712_not
g3563 not n715 ; n715_not
g3564 not n717 ; n717_not
g3565 not n719 ; n719_not
g3566 not n708 ; n708_not
g3567 not n720 ; n720_not
g3568 not n723 ; n723_not
g3569 not n725 ; n725_not
g3570 not n728 ; n728_not
g3571 not n730 ; n730_not
g3572 not n732 ; n732_not
g3573 not n735 ; n735_not
g3574 not n737 ; n737_not
g3575 not n740 ; n740_not
g3576 not n742 ; n742_not
g3577 not n744 ; n744_not
g3578 not n733 ; n733_not
g3579 not n745 ; n745_not
g3580 not n747 ; n747_not
g3581 not n750 ; n750_not
g3582 not n752 ; n752_not
g3583 not n755 ; n755_not
g3584 not n757 ; n757_not
g3585 not n759 ; n759_not
g3586 not n762 ; n762_not
g3587 not n764 ; n764_not
g3588 not n767 ; n767_not
g3589 not n769 ; n769_not
g3590 not n771 ; n771_not
g3591 not n760 ; n760_not
g3592 not n772 ; n772_not
g3593 not n775 ; n775_not
g3594 not n777 ; n777_not
g3595 not n780 ; n780_not
g3596 not n782 ; n782_not
g3597 not n784 ; n784_not
g3598 not n787 ; n787_not
g3599 not n789 ; n789_not
g3600 not n792 ; n792_not
g3601 not n794 ; n794_not
g3602 not n796 ; n796_not
g3603 not n785 ; n785_not
g3604 not n797 ; n797_not
g3605 not n799 ; n799_not
g3606 not n748 ; n748_not
g3607 not n800 ; n800_not
g3608 not n803 ; n803_not
g3609 not n805 ; n805_not
g3610 not n808 ; n808_not
g3611 not n810 ; n810_not
g3612 not n812 ; n812_not
g3613 not n815 ; n815_not
g3614 not n817 ; n817_not
g3615 not n820 ; n820_not
g3616 not n822 ; n822_not
g3617 not n824 ; n824_not
g3618 not n813 ; n813_not
g3619 not n825 ; n825_not
g3620 not n828 ; n828_not
g3621 not n830 ; n830_not
g3622 not n833 ; n833_not
g3623 not n835 ; n835_not
g3624 not n837 ; n837_not
g3625 not n840 ; n840_not
g3626 not n842 ; n842_not
g3627 not n845 ; n845_not
g3628 not n847 ; n847_not
g3629 not n849 ; n849_not
g3630 not n838 ; n838_not
g3631 not n850 ; n850_not
g3632 not n852 ; n852_not
g3633 not n855 ; n855_not
g3634 not n857 ; n857_not
g3635 not n860 ; n860_not
g3636 not n862 ; n862_not
g3637 not n864 ; n864_not
g3638 not n867 ; n867_not
g3639 not n869 ; n869_not
g3640 not n872 ; n872_not
g3641 not n874 ; n874_not
g3642 not n876 ; n876_not
g3643 not n865 ; n865_not
g3644 not n877 ; n877_not
g3645 not n880 ; n880_not
g3646 not n882 ; n882_not
g3647 not n885 ; n885_not
g3648 not n887 ; n887_not
g3649 not n889 ; n889_not
g3650 not n892 ; n892_not
g3651 not n894 ; n894_not
g3652 not n897 ; n897_not
g3653 not n899 ; n899_not
g3654 not n901 ; n901_not
g3655 not n890 ; n890_not
g3656 not n902 ; n902_not
g3657 not n904 ; n904_not
g3658 not n853 ; n853_not
g3659 not n905 ; n905_not
g3660 not n907 ; n907_not
g3661 not n910 ; n910_not
g3662 not n912 ; n912_not
g3663 not n915 ; n915_not
g3664 not n917 ; n917_not
g3665 not n919 ; n919_not
g3666 not n922 ; n922_not
g3667 not n924 ; n924_not
g3668 not n927 ; n927_not
g3669 not n929 ; n929_not
g3670 not n931 ; n931_not
g3671 not n920 ; n920_not
g3672 not n932 ; n932_not
g3673 not n935 ; n935_not
g3674 not n937 ; n937_not
g3675 not n940 ; n940_not
g3676 not n942 ; n942_not
g3677 not n944 ; n944_not
g3678 not n947 ; n947_not
g3679 not n949 ; n949_not
g3680 not n952 ; n952_not
g3681 not n954 ; n954_not
g3682 not n956 ; n956_not
g3683 not n945 ; n945_not
g3684 not n957 ; n957_not
g3685 not n959 ; n959_not
g3686 not n962 ; n962_not
g3687 not n964 ; n964_not
g3688 not n967 ; n967_not
g3689 not n969 ; n969_not
g3690 not n971 ; n971_not
g3691 not n974 ; n974_not
g3692 not n976 ; n976_not
g3693 not n979 ; n979_not
g3694 not n981 ; n981_not
g3695 not n983 ; n983_not
g3696 not n972 ; n972_not
g3697 not n984 ; n984_not
g3698 not n987 ; n987_not
g3699 not n989 ; n989_not
g3700 not n992 ; n992_not
g3701 not n994 ; n994_not
g3702 not n996 ; n996_not
g3703 not n999 ; n999_not
g3704 not n1001 ; n1001_not
g3705 not n1004 ; n1004_not
g3706 not n1006 ; n1006_not
g3707 not n1008 ; n1008_not
g3708 not n997 ; n997_not
g3709 not n1009 ; n1009_not
g3710 not n1011 ; n1011_not
g3711 not n960 ; n960_not
g3712 not n1012 ; n1012_not
g3713 not n1015 ; n1015_not
g3714 not n1017 ; n1017_not
g3715 not n1020 ; n1020_not
g3716 not n1022 ; n1022_not
g3717 not n1024 ; n1024_not
g3718 not n1027 ; n1027_not
g3719 not n1029 ; n1029_not
g3720 not n1032 ; n1032_not
g3721 not n1034 ; n1034_not
g3722 not n1036 ; n1036_not
g3723 not n1025 ; n1025_not
g3724 not n1037 ; n1037_not
g3725 not n1040 ; n1040_not
g3726 not n1042 ; n1042_not
g3727 not n1045 ; n1045_not
g3728 not n1047 ; n1047_not
g3729 not n1049 ; n1049_not
g3730 not n1052 ; n1052_not
g3731 not n1054 ; n1054_not
g3732 not n1057 ; n1057_not
g3733 not n1059 ; n1059_not
g3734 not n1061 ; n1061_not
g3735 not n1050 ; n1050_not
g3736 not n1062 ; n1062_not
g3737 not n1064 ; n1064_not
g3738 not n1067 ; n1067_not
g3739 not n1069 ; n1069_not
g3740 not n1072 ; n1072_not
g3741 not n1074 ; n1074_not
g3742 not n1076 ; n1076_not
g3743 not n1079 ; n1079_not
g3744 not n1081 ; n1081_not
g3745 not n1084 ; n1084_not
g3746 not n1086 ; n1086_not
g3747 not n1088 ; n1088_not
g3748 not n1077 ; n1077_not
g3749 not n1089 ; n1089_not
g3750 not n1092 ; n1092_not
g3751 not n1094 ; n1094_not
g3752 not n1097 ; n1097_not
g3753 not n1099 ; n1099_not
g3754 not n1101 ; n1101_not
g3755 not n1104 ; n1104_not
g3756 not n1106 ; n1106_not
g3757 not n1109 ; n1109_not
g3758 not n1111 ; n1111_not
g3759 not n1113 ; n1113_not
g3760 not n1102 ; n1102_not
g3761 not n1114 ; n1114_not
g3762 not n1116 ; n1116_not
g3763 not n1065 ; n1065_not
g3764 not n1117 ; n1117_not
g3765 not n1119 ; n1119_not
g3766 not n908 ; n908_not
g3767 not n1120 ; n1120_not
g3768 not n1122 ; n1122_not
g3769 not n1123 ; n1123_not
g3770 not n1125 ; n1125_not
g3771 not n1126 ; n1126_not
g3772 not n1128 ; n1128_not
g3773 not n1130 ; n1130_not
g3774 not n1131 ; n1131_not
g3775 not n1133 ; n1133_not
g3776 not n1134 ; n1134_not
g3777 not n1136 ; n1136_not
g3778 not n1129 ; n1129_not
g3779 not n1137 ; n1137_not
g3780 not n1139 ; n1139_not
g3781 not n1140 ; n1140_not
g3782 not n1142 ; n1142_not
g3783 not n1143 ; n1143_not
g3784 not n1145 ; n1145_not
g3785 not n1147 ; n1147_not
g3786 not n1148 ; n1148_not
g3787 not n1150 ; n1150_not
g3788 not n1151 ; n1151_not
g3789 not n1153 ; n1153_not
g3790 not n1146 ; n1146_not
g3791 not n1154 ; n1154_not
g3792 not n1156 ; n1156_not
g3793 not n1158 ; n1158_not
g3794 not n1159 ; n1159_not
g3795 not n1161 ; n1161_not
g3796 not n1162 ; n1162_not
g3797 not n1164 ; n1164_not
g3798 not n1166 ; n1166_not
g3799 not n1167 ; n1167_not
g3800 not n1169 ; n1169_not
g3801 not n1170 ; n1170_not
g3802 not n1172 ; n1172_not
g3803 not n1165 ; n1165_not
g3804 not n1173 ; n1173_not
g3805 not n1175 ; n1175_not
g3806 not n1176 ; n1176_not
g3807 not n1178 ; n1178_not
g3808 not n1179 ; n1179_not
g3809 not n1181 ; n1181_not
g3810 not n1183 ; n1183_not
g3811 not n1184 ; n1184_not
g3812 not n1186 ; n1186_not
g3813 not n1187 ; n1187_not
g3814 not n1189 ; n1189_not
g3815 not n1182 ; n1182_not
g3816 not n1190 ; n1190_not
g3817 not n1192 ; n1192_not
g3818 not n1157 ; n1157_not
g3819 not n1193 ; n1193_not
g3820 not n1195 ; n1195_not
g3821 not n1196 ; n1196_not
g3822 not n1198 ; n1198_not
g3823 not n1199 ; n1199_not
g3824 not n1201 ; n1201_not
g3825 not n1203 ; n1203_not
g3826 not n1204 ; n1204_not
g3827 not n1206 ; n1206_not
g3828 not n1207 ; n1207_not
g3829 not n1209 ; n1209_not
g3830 not n1202 ; n1202_not
g3831 not n1210 ; n1210_not
g3832 not n1212 ; n1212_not
g3833 not n1213 ; n1213_not
g3834 not n1215 ; n1215_not
g3835 not n1216 ; n1216_not
g3836 not n1218 ; n1218_not
g3837 not n1220 ; n1220_not
g3838 not n1221 ; n1221_not
g3839 not n1223 ; n1223_not
g3840 not n1224 ; n1224_not
g3841 not n1226 ; n1226_not
g3842 not n1219 ; n1219_not
g3843 not n1227 ; n1227_not
g3844 not n1229 ; n1229_not
g3845 not n1231 ; n1231_not
g3846 not n1232 ; n1232_not
g3847 not n1234 ; n1234_not
g3848 not n1235 ; n1235_not
g3849 not n1237 ; n1237_not
g3850 not n1239 ; n1239_not
g3851 not n1240 ; n1240_not
g3852 not n1242 ; n1242_not
g3853 not n1243 ; n1243_not
g3854 not n1245 ; n1245_not
g3855 not n1238 ; n1238_not
g3856 not n1246 ; n1246_not
g3857 not n1248 ; n1248_not
g3858 not n1249 ; n1249_not
g3859 not n1251 ; n1251_not
g3860 not n1252 ; n1252_not
g3861 not n1254 ; n1254_not
g3862 not n1256 ; n1256_not
g3863 not n1257 ; n1257_not
g3864 not n1259 ; n1259_not
g3865 not n1260 ; n1260_not
g3866 not n1262 ; n1262_not
g3867 not n1255 ; n1255_not
g3868 not n1263 ; n1263_not
g3869 not n1265 ; n1265_not
g3870 not n1230 ; n1230_not
g3871 not n1266 ; n1266_not
g3872 not n1268 ; n1268_not
g3873 not n1270 ; n1270_not
g3874 not n1271 ; n1271_not
g3875 not n1273 ; n1273_not
g3876 not n1274 ; n1274_not
g3877 not n1276 ; n1276_not
g3878 not n1278 ; n1278_not
g3879 not n1279 ; n1279_not
g3880 not n1281 ; n1281_not
g3881 not n1282 ; n1282_not
g3882 not n1284 ; n1284_not
g3883 not n1277 ; n1277_not
g3884 not n1285 ; n1285_not
g3885 not n1287 ; n1287_not
g3886 not n1288 ; n1288_not
g3887 not n1290 ; n1290_not
g3888 not n1291 ; n1291_not
g3889 not n1293 ; n1293_not
g3890 not n1295 ; n1295_not
g3891 not n1296 ; n1296_not
g3892 not n1298 ; n1298_not
g3893 not n1299 ; n1299_not
g3894 not n1301 ; n1301_not
g3895 not n1294 ; n1294_not
g3896 not n1302 ; n1302_not
g3897 not n1304 ; n1304_not
g3898 not n1306 ; n1306_not
g3899 not n1307 ; n1307_not
g3900 not n1309 ; n1309_not
g3901 not n1310 ; n1310_not
g3902 not n1312 ; n1312_not
g3903 not n1314 ; n1314_not
g3904 not n1315 ; n1315_not
g3905 not n1317 ; n1317_not
g3906 not n1318 ; n1318_not
g3907 not n1320 ; n1320_not
g3908 not n1313 ; n1313_not
g3909 not n1321 ; n1321_not
g3910 not n1323 ; n1323_not
g3911 not n1324 ; n1324_not
g3912 not n1326 ; n1326_not
g3913 not n1327 ; n1327_not
g3914 not n1329 ; n1329_not
g3915 not n1331 ; n1331_not
g3916 not n1332 ; n1332_not
g3917 not n1334 ; n1334_not
g3918 not n1335 ; n1335_not
g3919 not n1337 ; n1337_not
g3920 not n1330 ; n1330_not
g3921 not n1338 ; n1338_not
g3922 not n1340 ; n1340_not
g3923 not n1305 ; n1305_not
g3924 not n1341 ; n1341_not
g3925 not n1343 ; n1343_not
g3926 not n1344 ; n1344_not
g3927 not n1346 ; n1346_not
g3928 not n1347 ; n1347_not
g3929 not n1349 ; n1349_not
g3930 not n1351 ; n1351_not
g3931 not n1352 ; n1352_not
g3932 not n1354 ; n1354_not
g3933 not n1355 ; n1355_not
g3934 not n1357 ; n1357_not
g3935 not n1350 ; n1350_not
g3936 not n1358 ; n1358_not
g3937 not n1360 ; n1360_not
g3938 not n1361 ; n1361_not
g3939 not n1363 ; n1363_not
g3940 not n1364 ; n1364_not
g3941 not n1366 ; n1366_not
g3942 not n1368 ; n1368_not
g3943 not n1369 ; n1369_not
g3944 not n1371 ; n1371_not
g3945 not n1372 ; n1372_not
g3946 not n1374 ; n1374_not
g3947 not n1367 ; n1367_not
g3948 not n1375 ; n1375_not
g3949 not n1377 ; n1377_not
g3950 not n1379 ; n1379_not
g3951 not n1380 ; n1380_not
g3952 not n1382 ; n1382_not
g3953 not n1383 ; n1383_not
g3954 not n1385 ; n1385_not
g3955 not n1387 ; n1387_not
g3956 not n1388 ; n1388_not
g3957 not n1390 ; n1390_not
g3958 not n1391 ; n1391_not
g3959 not n1393 ; n1393_not
g3960 not n1386 ; n1386_not
g3961 not n1394 ; n1394_not
g3962 not n1396 ; n1396_not
g3963 not n1397 ; n1397_not
g3964 not n1399 ; n1399_not
g3965 not n1400 ; n1400_not
g3966 not n1402 ; n1402_not
g3967 not n1404 ; n1404_not
g3968 not n1405 ; n1405_not
g3969 not n1407 ; n1407_not
g3970 not n1408 ; n1408_not
g3971 not n1410 ; n1410_not
g3972 not n1403 ; n1403_not
g3973 not n1411 ; n1411_not
g3974 not n1413 ; n1413_not
g3975 not n1378 ; n1378_not
g3976 not n1414 ; n1414_not
g3977 not n1416 ; n1416_not
g3978 not n1269 ; n1269_not
g3979 not n1417 ; n1417_not
g3980 not n1419 ; n1419_not
g3981 not n1420 ; n1420_not
g3982 not n1422 ; n1422_not
g3983 not n1423 ; n1423_not
g3984 not n1425 ; n1425_not
g3985 not n1427 ; n1427_not
g3986 not n1428 ; n1428_not
g3987 not n1430 ; n1430_not
g3988 not n1431 ; n1431_not
g3989 not n1433 ; n1433_not
g3990 not n1426 ; n1426_not
g3991 not n1434 ; n1434_not
g3992 not n1436 ; n1436_not
g3993 not n1437 ; n1437_not
g3994 not n1439 ; n1439_not
g3995 not n1440 ; n1440_not
g3996 not n1442 ; n1442_not
g3997 not n1444 ; n1444_not
g3998 not n1445 ; n1445_not
g3999 not n1447 ; n1447_not
g4000 not n1448 ; n1448_not
g4001 not n1450 ; n1450_not
g4002 not n1443 ; n1443_not
g4003 not n1451 ; n1451_not
g4004 not n1453 ; n1453_not
g4005 not n1455 ; n1455_not
g4006 not n1456 ; n1456_not
g4007 not n1458 ; n1458_not
g4008 not n1459 ; n1459_not
g4009 not n1461 ; n1461_not
g4010 not n1463 ; n1463_not
g4011 not n1464 ; n1464_not
g4012 not n1466 ; n1466_not
g4013 not n1467 ; n1467_not
g4014 not n1469 ; n1469_not
g4015 not n1462 ; n1462_not
g4016 not n1470 ; n1470_not
g4017 not n1472 ; n1472_not
g4018 not n1473 ; n1473_not
g4019 not n1475 ; n1475_not
g4020 not n1476 ; n1476_not
g4021 not n1478 ; n1478_not
g4022 not n1480 ; n1480_not
g4023 not n1481 ; n1481_not
g4024 not n1483 ; n1483_not
g4025 not n1484 ; n1484_not
g4026 not n1486 ; n1486_not
g4027 not n1479 ; n1479_not
g4028 not n1487 ; n1487_not
g4029 not n1489 ; n1489_not
g4030 not n1454 ; n1454_not
g4031 not n1490 ; n1490_not
g4032 not n1492 ; n1492_not
g4033 not n1493 ; n1493_not
g4034 not n1495 ; n1495_not
g4035 not n1496 ; n1496_not
g4036 not n1498 ; n1498_not
g4037 not n1500 ; n1500_not
g4038 not n1501 ; n1501_not
g4039 not n1503 ; n1503_not
g4040 not n1504 ; n1504_not
g4041 not n1506 ; n1506_not
g4042 not n1499 ; n1499_not
g4043 not n1507 ; n1507_not
g4044 not n1509 ; n1509_not
g4045 not n1510 ; n1510_not
g4046 not n1512 ; n1512_not
g4047 not n1513 ; n1513_not
g4048 not n1515 ; n1515_not
g4049 not n1517 ; n1517_not
g4050 not n1518 ; n1518_not
g4051 not n1520 ; n1520_not
g4052 not n1521 ; n1521_not
g4053 not n1523 ; n1523_not
g4054 not n1516 ; n1516_not
g4055 not n1524 ; n1524_not
g4056 not n1526 ; n1526_not
g4057 not n1528 ; n1528_not
g4058 not n1529 ; n1529_not
g4059 not n1531 ; n1531_not
g4060 not n1532 ; n1532_not
g4061 not n1534 ; n1534_not
g4062 not n1536 ; n1536_not
g4063 not n1537 ; n1537_not
g4064 not n1539 ; n1539_not
g4065 not n1540 ; n1540_not
g4066 not n1542 ; n1542_not
g4067 not n1535 ; n1535_not
g4068 not n1543 ; n1543_not
g4069 not n1545 ; n1545_not
g4070 not n1546 ; n1546_not
g4071 not n1548 ; n1548_not
g4072 not n1549 ; n1549_not
g4073 not n1551 ; n1551_not
g4074 not n1553 ; n1553_not
g4075 not n1554 ; n1554_not
g4076 not n1556 ; n1556_not
g4077 not n1557 ; n1557_not
g4078 not n1559 ; n1559_not
g4079 not n1552 ; n1552_not
g4080 not n1560 ; n1560_not
g4081 not n1562 ; n1562_not
g4082 not n1527 ; n1527_not
g4083 not n1563 ; n1563_not
g4084 not n1565 ; n1565_not
g4085 not n1567 ; n1567_not
g4086 not n1568 ; n1568_not
g4087 not n1570 ; n1570_not
g4088 not n1571 ; n1571_not
g4089 not n1573 ; n1573_not
g4090 not n1575 ; n1575_not
g4091 not n1576 ; n1576_not
g4092 not n1578 ; n1578_not
g4093 not n1579 ; n1579_not
g4094 not n1581 ; n1581_not
g4095 not n1574 ; n1574_not
g4096 not n1582 ; n1582_not
g4097 not n1584 ; n1584_not
g4098 not n1585 ; n1585_not
g4099 not n1587 ; n1587_not
g4100 not n1588 ; n1588_not
g4101 not n1590 ; n1590_not
g4102 not n1592 ; n1592_not
g4103 not n1593 ; n1593_not
g4104 not n1595 ; n1595_not
g4105 not n1596 ; n1596_not
g4106 not n1598 ; n1598_not
g4107 not n1591 ; n1591_not
g4108 not n1599 ; n1599_not
g4109 not n1601 ; n1601_not
g4110 not n1603 ; n1603_not
g4111 not n1604 ; n1604_not
g4112 not n1606 ; n1606_not
g4113 not n1607 ; n1607_not
g4114 not n1609 ; n1609_not
g4115 not n1611 ; n1611_not
g4116 not n1612 ; n1612_not
g4117 not n1614 ; n1614_not
g4118 not n1615 ; n1615_not
g4119 not n1617 ; n1617_not
g4120 not n1610 ; n1610_not
g4121 not n1618 ; n1618_not
g4122 not n1620 ; n1620_not
g4123 not n1621 ; n1621_not
g4124 not n1623 ; n1623_not
g4125 not n1624 ; n1624_not
g4126 not n1626 ; n1626_not
g4127 not n1628 ; n1628_not
g4128 not n1629 ; n1629_not
g4129 not n1631 ; n1631_not
g4130 not n1632 ; n1632_not
g4131 not n1634 ; n1634_not
g4132 not n1627 ; n1627_not
g4133 not n1635 ; n1635_not
g4134 not n1637 ; n1637_not
g4135 not n1602 ; n1602_not
g4136 not n1638 ; n1638_not
g4137 not n1640 ; n1640_not
g4138 not n1641 ; n1641_not
g4139 not n1643 ; n1643_not
g4140 not n1644 ; n1644_not
g4141 not n1646 ; n1646_not
g4142 not n1648 ; n1648_not
g4143 not n1649 ; n1649_not
g4144 not n1651 ; n1651_not
g4145 not n1652 ; n1652_not
g4146 not n1654 ; n1654_not
g4147 not n1647 ; n1647_not
g4148 not n1655 ; n1655_not
g4149 not n1657 ; n1657_not
g4150 not n1658 ; n1658_not
g4151 not n1660 ; n1660_not
g4152 not n1661 ; n1661_not
g4153 not n1663 ; n1663_not
g4154 not n1665 ; n1665_not
g4155 not n1666 ; n1666_not
g4156 not n1668 ; n1668_not
g4157 not n1669 ; n1669_not
g4158 not n1671 ; n1671_not
g4159 not n1664 ; n1664_not
g4160 not n1672 ; n1672_not
g4161 not n1674 ; n1674_not
g4162 not n1676 ; n1676_not
g4163 not n1677 ; n1677_not
g4164 not n1679 ; n1679_not
g4165 not n1680 ; n1680_not
g4166 not n1682 ; n1682_not
g4167 not n1684 ; n1684_not
g4168 not n1685 ; n1685_not
g4169 not n1687 ; n1687_not
g4170 not n1688 ; n1688_not
g4171 not n1690 ; n1690_not
g4172 not n1683 ; n1683_not
g4173 not n1691 ; n1691_not
g4174 not n1693 ; n1693_not
g4175 not n1694 ; n1694_not
g4176 not n1696 ; n1696_not
g4177 not n1697 ; n1697_not
g4178 not n1699 ; n1699_not
g4179 not n1701 ; n1701_not
g4180 not n1702 ; n1702_not
g4181 not n1704 ; n1704_not
g4182 not n1705 ; n1705_not
g4183 not n1707 ; n1707_not
g4184 not n1700 ; n1700_not
g4185 not n1708 ; n1708_not
g4186 not n1710 ; n1710_not
g4187 not n1675 ; n1675_not
g4188 not n1711 ; n1711_not
g4189 not n1713 ; n1713_not
g4190 not n1566 ; n1566_not
g4191 not n1714 ; n1714_not
g4192 not n1716 ; n1716_not
g4193 not n1717 ; n1717_not
g4194 not n1719 ; n1719_not
g4195 not n1720 ; n1720_not
g4196 not n1722 ; n1722_not
g4197 not n1724 ; n1724_not
g4198 not n1725 ; n1725_not
g4199 not n1727 ; n1727_not
g4200 not n1728 ; n1728_not
g4201 not n1730 ; n1730_not
g4202 not n1723 ; n1723_not
g4203 not n1731 ; n1731_not
g4204 not n1733 ; n1733_not
g4205 not n1734 ; n1734_not
g4206 not n1736 ; n1736_not
g4207 not n1737 ; n1737_not
g4208 not n1739 ; n1739_not
g4209 not n1741 ; n1741_not
g4210 not n1742 ; n1742_not
g4211 not n1744 ; n1744_not
g4212 not n1745 ; n1745_not
g4213 not n1747 ; n1747_not
g4214 not n1740 ; n1740_not
g4215 not n1748 ; n1748_not
g4216 not n1750 ; n1750_not
g4217 not n1752 ; n1752_not
g4218 not n1753 ; n1753_not
g4219 not n1755 ; n1755_not
g4220 not n1756 ; n1756_not
g4221 not n1758 ; n1758_not
g4222 not n1760 ; n1760_not
g4223 not n1761 ; n1761_not
g4224 not n1763 ; n1763_not
g4225 not n1764 ; n1764_not
g4226 not n1766 ; n1766_not
g4227 not n1759 ; n1759_not
g4228 not n1767 ; n1767_not
g4229 not n1769 ; n1769_not
g4230 not n1770 ; n1770_not
g4231 not n1772 ; n1772_not
g4232 not n1773 ; n1773_not
g4233 not n1775 ; n1775_not
g4234 not n1777 ; n1777_not
g4235 not n1778 ; n1778_not
g4236 not n1780 ; n1780_not
g4237 not n1781 ; n1781_not
g4238 not n1783 ; n1783_not
g4239 not n1776 ; n1776_not
g4240 not n1784 ; n1784_not
g4241 not n1786 ; n1786_not
g4242 not n1751 ; n1751_not
g4243 not n1787 ; n1787_not
g4244 not n1789 ; n1789_not
g4245 not n1790 ; n1790_not
g4246 not n1792 ; n1792_not
g4247 not n1793 ; n1793_not
g4248 not n1795 ; n1795_not
g4249 not n1797 ; n1797_not
g4250 not n1798 ; n1798_not
g4251 not n1800 ; n1800_not
g4252 not n1801 ; n1801_not
g4253 not n1803 ; n1803_not
g4254 not n1796 ; n1796_not
g4255 not n1804 ; n1804_not
g4256 not n1806 ; n1806_not
g4257 not n1807 ; n1807_not
g4258 not n1809 ; n1809_not
g4259 not n1810 ; n1810_not
g4260 not n1812 ; n1812_not
g4261 not n1814 ; n1814_not
g4262 not n1815 ; n1815_not
g4263 not n1817 ; n1817_not
g4264 not n1818 ; n1818_not
g4265 not n1820 ; n1820_not
g4266 not n1813 ; n1813_not
g4267 not n1821 ; n1821_not
g4268 not n1823 ; n1823_not
g4269 not n1825 ; n1825_not
g4270 not n1826 ; n1826_not
g4271 not n1828 ; n1828_not
g4272 not n1829 ; n1829_not
g4273 not n1831 ; n1831_not
g4274 not n1833 ; n1833_not
g4275 not n1834 ; n1834_not
g4276 not n1836 ; n1836_not
g4277 not n1837 ; n1837_not
g4278 not n1839 ; n1839_not
g4279 not n1832 ; n1832_not
g4280 not n1840 ; n1840_not
g4281 not n1842 ; n1842_not
g4282 not n1843 ; n1843_not
g4283 not n1845 ; n1845_not
g4284 not n1846 ; n1846_not
g4285 not n1848 ; n1848_not
g4286 not n1850 ; n1850_not
g4287 not n1851 ; n1851_not
g4288 not n1853 ; n1853_not
g4289 not n1854 ; n1854_not
g4290 not n1856 ; n1856_not
g4291 not n1849 ; n1849_not
g4292 not n1857 ; n1857_not
g4293 not n1859 ; n1859_not
g4294 not n1824 ; n1824_not
g4295 not n1860 ; n1860_not
g4296 not n1862 ; n1862_not
g4297 not n1863 ; n1863_not
g4298 not n1865 ; n1865_not
g4299 not n1866 ; n1866_not
g4300 not n1868 ; n1868_not
g4301 not n1870 ; n1870_not
g4302 not n1871 ; n1871_not
g4303 not n1873 ; n1873_not
g4304 not n1874 ; n1874_not
g4305 not n1876 ; n1876_not
g4306 not n1869 ; n1869_not
g4307 not n1877 ; n1877_not
g4308 not n1879 ; n1879_not
g4309 not n1880 ; n1880_not
g4310 not n1882 ; n1882_not
g4311 not n1883 ; n1883_not
g4312 not n1885 ; n1885_not
g4313 not n1887 ; n1887_not
g4314 not n1888 ; n1888_not
g4315 not n1890 ; n1890_not
g4316 not n1891 ; n1891_not
g4317 not n1893 ; n1893_not
g4318 not n1886 ; n1886_not
g4319 not n1894 ; n1894_not
g4320 not n1896 ; n1896_not
g4321 not n1898 ; n1898_not
g4322 not n1899 ; n1899_not
g4323 not n1901 ; n1901_not
g4324 not n1902 ; n1902_not
g4325 not n1904 ; n1904_not
g4326 not n1906 ; n1906_not
g4327 not n1907 ; n1907_not
g4328 not n1909 ; n1909_not
g4329 not n1910 ; n1910_not
g4330 not n1912 ; n1912_not
g4331 not n1905 ; n1905_not
g4332 not n1913 ; n1913_not
g4333 not n1915 ; n1915_not
g4334 not n1916 ; n1916_not
g4335 not n1918 ; n1918_not
g4336 not n1919 ; n1919_not
g4337 not n1921 ; n1921_not
g4338 not n1923 ; n1923_not
g4339 not n1924 ; n1924_not
g4340 not n1926 ; n1926_not
g4341 not n1927 ; n1927_not
g4342 not n1929 ; n1929_not
g4343 not n1922 ; n1922_not
g4344 not n1930 ; n1930_not
g4345 not n1932 ; n1932_not
g4346 not n1897 ; n1897_not
g4347 not n1933 ; n1933_not
g4348 not n1935 ; n1935_not
g4349 not n1936 ; n1936_not
g4350 not n1938 ; n1938_not
g4351 not n1939 ; n1939_not
g4352 not n1941 ; n1941_not
g4353 not n1943 ; n1943_not
g4354 not n1944 ; n1944_not
g4355 not n1946 ; n1946_not
g4356 not n1947 ; n1947_not
g4357 not n1949 ; n1949_not
g4358 not n1942 ; n1942_not
g4359 not n1950 ; n1950_not
g4360 not n1952 ; n1952_not
g4361 not n1953 ; n1953_not
g4362 not n1955 ; n1955_not
g4363 not n1956 ; n1956_not
g4364 not n1958 ; n1958_not
g4365 not n1960 ; n1960_not
g4366 not n1961 ; n1961_not
g4367 not n1963 ; n1963_not
g4368 not n1964 ; n1964_not
g4369 not n1966 ; n1966_not
g4370 not n1959 ; n1959_not
g4371 not n1967 ; n1967_not
g4372 not n1969 ; n1969_not
g4373 not n1971 ; n1971_not
g4374 not n1972 ; n1972_not
g4375 not n1974 ; n1974_not
g4376 not n1975 ; n1975_not
g4377 not n1977 ; n1977_not
g4378 not n1979 ; n1979_not
g4379 not n1980 ; n1980_not
g4380 not n1982 ; n1982_not
g4381 not n1983 ; n1983_not
g4382 not n1985 ; n1985_not
g4383 not n1978 ; n1978_not
g4384 not n1986 ; n1986_not
g4385 not n1988 ; n1988_not
g4386 not n1989 ; n1989_not
g4387 not n1991 ; n1991_not
g4388 not n1992 ; n1992_not
g4389 not n1994 ; n1994_not
g4390 not n1996 ; n1996_not
g4391 not n1997 ; n1997_not
g4392 not n1999 ; n1999_not
g4393 not n2000 ; n2000_not
g4394 not n2002 ; n2002_not
g4395 not n1995 ; n1995_not
g4396 not n2003 ; n2003_not
g4397 not n2005 ; n2005_not
g4398 not n1970 ; n1970_not
g4399 not n2006 ; n2006_not
g4400 not n2008 ; n2008_not
g4401 not n2009 ; n2009_not
g4402 not n2011 ; n2011_not
g4403 not n2012 ; n2012_not
g4404 not n2014 ; n2014_not
g4405 not n2016 ; n2016_not
g4406 not n2017 ; n2017_not
g4407 not n2019 ; n2019_not
g4408 not n2020 ; n2020_not
g4409 not n2022 ; n2022_not
g4410 not n2015 ; n2015_not
g4411 not n2023 ; n2023_not
g4412 not n2025 ; n2025_not
g4413 not n2026 ; n2026_not
g4414 not n2028 ; n2028_not
g4415 not n2029 ; n2029_not
g4416 not n2031 ; n2031_not
g4417 not n2033 ; n2033_not
g4418 not n2034 ; n2034_not
g4419 not n2036 ; n2036_not
g4420 not n2037 ; n2037_not
g4421 not n2039 ; n2039_not
g4422 not n2032 ; n2032_not
g4423 not n2040 ; n2040_not
g4424 not n2042 ; n2042_not
g4425 not n2044 ; n2044_not
g4426 not n2045 ; n2045_not
g4427 not n2047 ; n2047_not
g4428 not n2048 ; n2048_not
g4429 not n2050 ; n2050_not
g4430 not n2052 ; n2052_not
g4431 not n2053 ; n2053_not
g4432 not n2055 ; n2055_not
g4433 not n2056 ; n2056_not
g4434 not n2058 ; n2058_not
g4435 not n2051 ; n2051_not
g4436 not n2059 ; n2059_not
g4437 not n2061 ; n2061_not
g4438 not n2062 ; n2062_not
g4439 not n2064 ; n2064_not
g4440 not n2065 ; n2065_not
g4441 not n2067 ; n2067_not
g4442 not n2069 ; n2069_not
g4443 not n2070 ; n2070_not
g4444 not n2072 ; n2072_not
g4445 not n2073 ; n2073_not
g4446 not n2075 ; n2075_not
g4447 not n2068 ; n2068_not
g4448 not n2076 ; n2076_not
g4449 not n2078 ; n2078_not
g4450 not n2043 ; n2043_not
g4451 not n2079 ; n2079_not
g4452 not n2081 ; n2081_not
g4453 not n2082 ; n2082_not
g4454 not n2084 ; n2084_not
g4455 not n2085 ; n2085_not
g4456 not n2087 ; n2087_not
g4457 not n2089 ; n2089_not
g4458 not n2090 ; n2090_not
g4459 not n2092 ; n2092_not
g4460 not n2093 ; n2093_not
g4461 not n2095 ; n2095_not
g4462 not n2088 ; n2088_not
g4463 not n2096 ; n2096_not
g4464 not n2098 ; n2098_not
g4465 not n2099 ; n2099_not
g4466 not n2101 ; n2101_not
g4467 not n2102 ; n2102_not
g4468 not n2104 ; n2104_not
g4469 not n2106 ; n2106_not
g4470 not n2107 ; n2107_not
g4471 not n2109 ; n2109_not
g4472 not n2110 ; n2110_not
g4473 not n2112 ; n2112_not
g4474 not n2105 ; n2105_not
g4475 not n2113 ; n2113_not
g4476 not n2115 ; n2115_not
g4477 not n2117 ; n2117_not
g4478 not n2118 ; n2118_not
g4479 not n2120 ; n2120_not
g4480 not n2121 ; n2121_not
g4481 not n2123 ; n2123_not
g4482 not n2125 ; n2125_not
g4483 not n2126 ; n2126_not
g4484 not n2128 ; n2128_not
g4485 not n2129 ; n2129_not
g4486 not n2131 ; n2131_not
g4487 not n2124 ; n2124_not
g4488 not n2132 ; n2132_not
g4489 not n2134 ; n2134_not
g4490 not n2135 ; n2135_not
g4491 not n2137 ; n2137_not
g4492 not n2138 ; n2138_not
g4493 not n2140 ; n2140_not
g4494 not n2142 ; n2142_not
g4495 not n2143 ; n2143_not
g4496 not n2145 ; n2145_not
g4497 not n2146 ; n2146_not
g4498 not n2148 ; n2148_not
g4499 not n2141 ; n2141_not
g4500 not n2149 ; n2149_not
g4501 not n2151 ; n2151_not
g4502 not n2116 ; n2116_not
g4503 not n2152 ; n2152_not
g4504 not n2154 ; n2154_not
g4505 not n2155 ; n2155_not
g4506 not n2157 ; n2157_not
g4507 not n2158 ; n2158_not
g4508 not n2160 ; n2160_not
g4509 not n2162 ; n2162_not
g4510 not n2163 ; n2163_not
g4511 not n2165 ; n2165_not
g4512 not n2166 ; n2166_not
g4513 not n2168 ; n2168_not
g4514 not n2161 ; n2161_not
g4515 not n2169 ; n2169_not
g4516 not n2171 ; n2171_not
g4517 not n2172 ; n2172_not
g4518 not n2174 ; n2174_not
g4519 not n2175 ; n2175_not
g4520 not n2177 ; n2177_not
g4521 not n2179 ; n2179_not
g4522 not n2180 ; n2180_not
g4523 not n2182 ; n2182_not
g4524 not n2183 ; n2183_not
g4525 not n2185 ; n2185_not
g4526 not n2178 ; n2178_not
g4527 not n2186 ; n2186_not
g4528 not n2188 ; n2188_not
g4529 not n2190 ; n2190_not
g4530 not n2191 ; n2191_not
g4531 not n2193 ; n2193_not
g4532 not n2194 ; n2194_not
g4533 not n2196 ; n2196_not
g4534 not n2198 ; n2198_not
g4535 not n2199 ; n2199_not
g4536 not n2201 ; n2201_not
g4537 not n2202 ; n2202_not
g4538 not n2204 ; n2204_not
g4539 not n2197 ; n2197_not
g4540 not n2205 ; n2205_not
g4541 not n2207 ; n2207_not
g4542 not n2208 ; n2208_not
g4543 not n2210 ; n2210_not
g4544 not n2211 ; n2211_not
g4545 not n2213 ; n2213_not
g4546 not n2215 ; n2215_not
g4547 not n2216 ; n2216_not
g4548 not n2218 ; n2218_not
g4549 not n2219 ; n2219_not
g4550 not n2221 ; n2221_not
g4551 not n2214 ; n2214_not
g4552 not n2222 ; n2222_not
g4553 not n2224 ; n2224_not
g4554 not n2189 ; n2189_not
g4555 not n2225 ; n2225_not
g4556 not n2227 ; n2227_not
g4557 not n2228 ; n2228_not
g4558 not n2230 ; n2230_not
g4559 not n2231 ; n2231_not
g4560 not n2233 ; n2233_not
g4561 not n2235 ; n2235_not
g4562 not n2236 ; n2236_not
g4563 not n2238 ; n2238_not
g4564 not n2239 ; n2239_not
g4565 not n2241 ; n2241_not
g4566 not n2234 ; n2234_not
g4567 not n2242 ; n2242_not
g4568 not n2244 ; n2244_not
g4569 not n2245 ; n2245_not
g4570 not n2247 ; n2247_not
g4571 not n2248 ; n2248_not
g4572 not n2250 ; n2250_not
g4573 not n2252 ; n2252_not
g4574 not n2253 ; n2253_not
g4575 not n2255 ; n2255_not
g4576 not n2256 ; n2256_not
g4577 not n2258 ; n2258_not
g4578 not n2251 ; n2251_not
g4579 not n2259 ; n2259_not
g4580 not n2261 ; n2261_not
g4581 not n2263 ; n2263_not
g4582 not n2264 ; n2264_not
g4583 not n2266 ; n2266_not
g4584 not n2267 ; n2267_not
g4585 not n2269 ; n2269_not
g4586 not n2271 ; n2271_not
g4587 not n2272 ; n2272_not
g4588 not n2274 ; n2274_not
g4589 not n2275 ; n2275_not
g4590 not n2277 ; n2277_not
g4591 not n2270 ; n2270_not
g4592 not n2278 ; n2278_not
g4593 not n2280 ; n2280_not
g4594 not n2281 ; n2281_not
g4595 not n2283 ; n2283_not
g4596 not n2284 ; n2284_not
g4597 not n2286 ; n2286_not
g4598 not n2288 ; n2288_not
g4599 not n2289 ; n2289_not
g4600 not n2291 ; n2291_not
g4601 not n2292 ; n2292_not
g4602 not n2294 ; n2294_not
g4603 not n2287 ; n2287_not
g4604 not n2295 ; n2295_not
g4605 not n2297 ; n2297_not
g4606 not n2262 ; n2262_not
g4607 not n2298 ; n2298_not
g4608 not n2300 ; n2300_not
g4609 not n2301 ; n2301_not
g4610 not n2303 ; n2303_not
g4611 not n2304 ; n2304_not
g4612 not n2306 ; n2306_not
g4613 not n2308 ; n2308_not
g4614 not n2309 ; n2309_not
g4615 not n2311 ; n2311_not
g4616 not n2312 ; n2312_not
g4617 not n2314 ; n2314_not
g4618 not n2307 ; n2307_not
g4619 not n2315 ; n2315_not
g4620 not n2317 ; n2317_not
g4621 not n2318 ; n2318_not
g4622 not n2320 ; n2320_not
g4623 not n2321 ; n2321_not
g4624 not n2323 ; n2323_not
g4625 not n2325 ; n2325_not
g4626 not n2326 ; n2326_not
g4627 not n2328 ; n2328_not
g4628 not n2329 ; n2329_not
g4629 not n2331 ; n2331_not
g4630 not n2324 ; n2324_not
g4631 not n2332 ; n2332_not
g4632 not n2334 ; n2334_not
g4633 not n2336 ; n2336_not
g4634 not n2337 ; n2337_not
g4635 not n2339 ; n2339_not
g4636 not n2340 ; n2340_not
g4637 not n2342 ; n2342_not
g4638 not n2344 ; n2344_not
g4639 not n2345 ; n2345_not
g4640 not n2347 ; n2347_not
g4641 not n2348 ; n2348_not
g4642 not n2350 ; n2350_not
g4643 not n2343 ; n2343_not
g4644 not n2351 ; n2351_not
g4645 not n2353 ; n2353_not
g4646 not n2354 ; n2354_not
g4647 not n2356 ; n2356_not
g4648 not n2357 ; n2357_not
g4649 not n2359 ; n2359_not
g4650 not n2361 ; n2361_not
g4651 not n2362 ; n2362_not
g4652 not n2364 ; n2364_not
g4653 not n2365 ; n2365_not
g4654 not n2367 ; n2367_not
g4655 not n2360 ; n2360_not
g4656 not n2368 ; n2368_not
g4657 not n2370 ; n2370_not
g4658 not n2335 ; n2335_not
g4659 not n2371 ; n2371_not
g4660 not n2373 ; n2373_not
g4661 not n2374 ; n2374_not
g4662 not n2376 ; n2376_not
g4663 not n2377 ; n2377_not
g4664 not n2379 ; n2379_not
g4665 not n2381 ; n2381_not
g4666 not n2382 ; n2382_not
g4667 not n2384 ; n2384_not
g4668 not n2385 ; n2385_not
g4669 not n2387 ; n2387_not
g4670 not n2380 ; n2380_not
g4671 not n2388 ; n2388_not
g4672 not n2390 ; n2390_not
g4673 not n2391 ; n2391_not
g4674 not n2393 ; n2393_not
g4675 not n2394 ; n2394_not
g4676 not n2396 ; n2396_not
g4677 not n2398 ; n2398_not
g4678 not n2399 ; n2399_not
g4679 not n2401 ; n2401_not
g4680 not n2402 ; n2402_not
g4681 not n2404 ; n2404_not
g4682 not n2397 ; n2397_not
g4683 not n2405 ; n2405_not
g4684 not n2407 ; n2407_not
g4685 not n2409 ; n2409_not
g4686 not n2410 ; n2410_not
g4687 not n2412 ; n2412_not
g4688 not n2413 ; n2413_not
g4689 not n2415 ; n2415_not
g4690 not n2417 ; n2417_not
g4691 not n2418 ; n2418_not
g4692 not n2420 ; n2420_not
g4693 not n2421 ; n2421_not
g4694 not n2423 ; n2423_not
g4695 not n2416 ; n2416_not
g4696 not n2424 ; n2424_not
g4697 not n2426 ; n2426_not
g4698 not n2427 ; n2427_not
g4699 not n2429 ; n2429_not
g4700 not n2430 ; n2430_not
g4701 not n2432 ; n2432_not
g4702 not n2434 ; n2434_not
g4703 not n2435 ; n2435_not
g4704 not n2437 ; n2437_not
g4705 not n2438 ; n2438_not
g4706 not n2440 ; n2440_not
g4707 not n2433 ; n2433_not
g4708 not n2441 ; n2441_not
g4709 not n2443 ; n2443_not
g4710 not n2408 ; n2408_not
g4711 not n2444 ; n2444_not
g4712 not n2446 ; n2446_not
g4713 not n2447 ; n2447_not
g4714 not n2449 ; n2449_not
g4715 not n2450 ; n2450_not
g4716 not n2452 ; n2452_not
g4717 not n2454 ; n2454_not
g4718 not n2455 ; n2455_not
g4719 not n2457 ; n2457_not
g4720 not n2458 ; n2458_not
g4721 not n2460 ; n2460_not
g4722 not n2453 ; n2453_not
g4723 not n2461 ; n2461_not
g4724 not n2463 ; n2463_not
g4725 not n2464 ; n2464_not
g4726 not n2466 ; n2466_not
g4727 not n2467 ; n2467_not
g4728 not n2469 ; n2469_not
g4729 not n2471 ; n2471_not
g4730 not n2472 ; n2472_not
g4731 not n2474 ; n2474_not
g4732 not n2475 ; n2475_not
g4733 not n2477 ; n2477_not
g4734 not n2470 ; n2470_not
g4735 not n2478 ; n2478_not
g4736 not n2480 ; n2480_not
g4737 not n2482 ; n2482_not
g4738 not n2483 ; n2483_not
g4739 not n2485 ; n2485_not
g4740 not n2486 ; n2486_not
g4741 not n2488 ; n2488_not
g4742 not n2490 ; n2490_not
g4743 not n2491 ; n2491_not
g4744 not n2493 ; n2493_not
g4745 not n2494 ; n2494_not
g4746 not n2496 ; n2496_not
g4747 not n2489 ; n2489_not
g4748 not n2497 ; n2497_not
g4749 not n2499 ; n2499_not
g4750 not n2500 ; n2500_not
g4751 not n2502 ; n2502_not
g4752 not n2503 ; n2503_not
g4753 not n2505 ; n2505_not
g4754 not n2507 ; n2507_not
g4755 not n2508 ; n2508_not
g4756 not n2510 ; n2510_not
g4757 not n2511 ; n2511_not
g4758 not n2513 ; n2513_not
g4759 not n2506 ; n2506_not
g4760 not n2514 ; n2514_not
g4761 not n2516 ; n2516_not
g4762 not n2481 ; n2481_not
g4763 not n2517 ; n2517_not
g4764 not n2519 ; n2519_not
g4765 not n2520 ; n2520_not
g4766 not n2522 ; n2522_not
g4767 not n2523 ; n2523_not
g4768 not n2525 ; n2525_not
g4769 not n2527 ; n2527_not
g4770 not n2528 ; n2528_not
g4771 not n2530 ; n2530_not
g4772 not n2531 ; n2531_not
g4773 not n2533 ; n2533_not
g4774 not n2526 ; n2526_not
g4775 not n2534 ; n2534_not
g4776 not n2536 ; n2536_not
g4777 not n2537 ; n2537_not
g4778 not n2539 ; n2539_not
g4779 not n2540 ; n2540_not
g4780 not n2542 ; n2542_not
g4781 not n2544 ; n2544_not
g4782 not n2545 ; n2545_not
g4783 not n2547 ; n2547_not
g4784 not n2548 ; n2548_not
g4785 not n2550 ; n2550_not
g4786 not n2543 ; n2543_not
g4787 not n2551 ; n2551_not
g4788 not n2553 ; n2553_not
g4789 not n2555 ; n2555_not
g4790 not n2556 ; n2556_not
g4791 not n2558 ; n2558_not
g4792 not n2559 ; n2559_not
g4793 not n2561 ; n2561_not
g4794 not n2563 ; n2563_not
g4795 not n2564 ; n2564_not
g4796 not n2566 ; n2566_not
g4797 not n2567 ; n2567_not
g4798 not n2569 ; n2569_not
g4799 not n2562 ; n2562_not
g4800 not n2570 ; n2570_not
g4801 not n2572 ; n2572_not
g4802 not n2573 ; n2573_not
g4803 not n2575 ; n2575_not
g4804 not n2576 ; n2576_not
g4805 not n2578 ; n2578_not
g4806 not n2580 ; n2580_not
g4807 not n2581 ; n2581_not
g4808 not n2583 ; n2583_not
g4809 not n2584 ; n2584_not
g4810 not n2586 ; n2586_not
g4811 not n2579 ; n2579_not
g4812 not n2587 ; n2587_not
g4813 not n2589 ; n2589_not
g4814 not n2554 ; n2554_not
g4815 not n2590 ; n2590_not
g4816 not n2592 ; n2592_not
g4817 not n2593 ; n2593_not
g4818 not n2595 ; n2595_not
g4819 not n2596 ; n2596_not
g4820 not n2598 ; n2598_not
g4821 not n2600 ; n2600_not
g4822 not n2601 ; n2601_not
g4823 not n2603 ; n2603_not
g4824 not n2604 ; n2604_not
g4825 not n2606 ; n2606_not
g4826 not n2599 ; n2599_not
g4827 not n2607 ; n2607_not
g4828 not n2609 ; n2609_not
g4829 not n2610 ; n2610_not
g4830 not n2612 ; n2612_not
g4831 not n2613 ; n2613_not
g4832 not n2615 ; n2615_not
g4833 not n2617 ; n2617_not
g4834 not n2618 ; n2618_not
g4835 not n2620 ; n2620_not
g4836 not n2621 ; n2621_not
g4837 not n2623 ; n2623_not
g4838 not n2616 ; n2616_not
g4839 not n2624 ; n2624_not
g4840 not n2626 ; n2626_not
g4841 not n2627 ; n2627_not
g4842 not n2629 ; n2629_not
g4843 not n2630 ; n2630_not
g4844 not n2632 ; n2632_not
g4845 not n2634 ; n2634_not
g4846 not n2635 ; n2635_not
g4847 not n2637 ; n2637_not
g4848 not n2638 ; n2638_not
g4849 not n2640 ; n2640_not
g4850 not n2633 ; n2633_not
g4851 not n2641 ; n2641_not
g4852 not n2643 ; n2643_not
g4853 not n2644 ; n2644_not
g4854 not n2646 ; n2646_not
g4855 not n2647 ; n2647_not
g4856 not n2649 ; n2649_not
g4857 not n2651 ; n2651_not
g4858 not n2652 ; n2652_not
g4859 not n2654 ; n2654_not
g4860 not n2655 ; n2655_not
g4861 not n2657 ; n2657_not
g4862 not n2650 ; n2650_not
g4863 not n2658 ; n2658_not
g4864 not n2660 ; n2660_not
g4865 not n2661 ; n2661_not
g4866 not n2663 ; n2663_not
g4867 not n2664 ; n2664_not
g4868 not n2666 ; n2666_not
g4869 not n2668 ; n2668_not
g4870 not n2669 ; n2669_not
g4871 not n2671 ; n2671_not
g4872 not n2672 ; n2672_not
g4873 not n2674 ; n2674_not
g4874 not n2667 ; n2667_not
g4875 not n2675 ; n2675_not
g4876 not n2677 ; n2677_not
g4877 not n2678 ; n2678_not
g4878 not n2680 ; n2680_not
g4879 not n2681 ; n2681_not
g4880 not n2683 ; n2683_not
g4881 not n2685 ; n2685_not
g4882 not n2686 ; n2686_not
g4883 not n2688 ; n2688_not
g4884 not n2689 ; n2689_not
g4885 not n2691 ; n2691_not
g4886 not n2684 ; n2684_not
g4887 not n2692 ; n2692_not
g4888 not n2694 ; n2694_not
g4889 not n2695 ; n2695_not
g4890 not n2697 ; n2697_not
g4891 not n2698 ; n2698_not
g4892 not n2700 ; n2700_not
g4893 not n2702 ; n2702_not
g4894 not n2703 ; n2703_not
g4895 not n2705 ; n2705_not
g4896 not n2706 ; n2706_not
g4897 not n2708 ; n2708_not
g4898 not n2701 ; n2701_not
g4899 not n2709 ; n2709_not
g4900 not n2711 ; n2711_not
g4901 not n2712 ; n2712_not
g4902 not n2714 ; n2714_not
g4903 not n2715 ; n2715_not
g4904 not n2717 ; n2717_not
g4905 not n2719 ; n2719_not
g4906 not n2720 ; n2720_not
g4907 not n2722 ; n2722_not
g4908 not n2723 ; n2723_not
g4909 not n2725 ; n2725_not
g4910 not n2718 ; n2718_not
g4911 not n2726 ; n2726_not
g4912 not n2728 ; n2728_not
g4913 not n2729 ; n2729_not
g4914 not n2731 ; n2731_not
g4915 not n2732 ; n2732_not
g4916 not n2734 ; n2734_not
g4917 not n2736 ; n2736_not
g4918 not n2737 ; n2737_not
g4919 not n2739 ; n2739_not
g4920 not n2740 ; n2740_not
g4921 not n2742 ; n2742_not
g4922 not n2735 ; n2735_not
g4923 not n2743 ; n2743_not
g4924 not n2745 ; n2745_not
g4925 not n2746 ; n2746_not
g4926 not n2748 ; n2748_not
g4927 not n2749 ; n2749_not
g4928 not n2751 ; n2751_not
g4929 not n2753 ; n2753_not
g4930 not n2754 ; n2754_not
g4931 not n2756 ; n2756_not
g4932 not n2757 ; n2757_not
g4933 not n2759 ; n2759_not
g4934 not n2752 ; n2752_not
g4935 not n2760 ; n2760_not
g4936 not n2762 ; n2762_not
g4937 not n2763 ; n2763_not
g4938 not n2765 ; n2765_not
g4939 not n2766 ; n2766_not
g4940 not n2768 ; n2768_not
g4941 not n2770 ; n2770_not
g4942 not n2771 ; n2771_not
g4943 not n2773 ; n2773_not
g4944 not n2774 ; n2774_not
g4945 not n2776 ; n2776_not
g4946 not n2769 ; n2769_not
g4947 not n2777 ; n2777_not
g4948 not n2779 ; n2779_not
g4949 not n2780 ; n2780_not
g4950 not n2782 ; n2782_not
g4951 not n2783 ; n2783_not
g4952 not n2785 ; n2785_not
g4953 not n2787 ; n2787_not
g4954 not n2788 ; n2788_not
g4955 not n2790 ; n2790_not
g4956 not n2791 ; n2791_not
g4957 not n2793 ; n2793_not
g4958 not n2786 ; n2786_not
g4959 not n2794 ; n2794_not
g4960 not n2796 ; n2796_not
g4961 not n2797 ; n2797_not
g4962 not n2799 ; n2799_not
g4963 not n2800 ; n2800_not
g4964 not n2802 ; n2802_not
g4965 not n2804 ; n2804_not
g4966 not n2805 ; n2805_not
g4967 not n2807 ; n2807_not
g4968 not n2808 ; n2808_not
g4969 not n2810 ; n2810_not
g4970 not n2803 ; n2803_not
g4971 not n2811 ; n2811_not
g4972 not n2813 ; n2813_not
g4973 not n2814 ; n2814_not
g4974 not n2816 ; n2816_not
g4975 not n2817 ; n2817_not
g4976 not n2819 ; n2819_not
g4977 not n2821 ; n2821_not
g4978 not n2822 ; n2822_not
g4979 not n2824 ; n2824_not
g4980 not n2825 ; n2825_not
g4981 not n2827 ; n2827_not
g4982 not n2820 ; n2820_not
g4983 not n2828 ; n2828_not
g4984 not n2830 ; n2830_not
g4985 not n2831 ; n2831_not
g4986 not n2833 ; n2833_not
g4987 not n2834 ; n2834_not
g4988 not n2836 ; n2836_not
g4989 not n2838 ; n2838_not
g4990 not n2839 ; n2839_not
g4991 not n2841 ; n2841_not
g4992 not n2842 ; n2842_not
g4993 not n2844 ; n2844_not
g4994 not n2837 ; n2837_not
g4995 not n2845 ; n2845_not
g4996 not n2847 ; n2847_not
g4997 not n2848 ; n2848_not
g4998 not n2850 ; n2850_not
g4999 not n2851 ; n2851_not
g5000 not n2853 ; n2853_not
g5001 not n2855 ; n2855_not
g5002 not n2856 ; n2856_not
g5003 not n2858 ; n2858_not
g5004 not n2859 ; n2859_not
g5005 not n2861 ; n2861_not
g5006 not n2854 ; n2854_not
g5007 not n2862 ; n2862_not
g5008 not n2864 ; n2864_not
g5009 not n2865 ; n2865_not
g5010 not n2867 ; n2867_not
g5011 not n2868 ; n2868_not
g5012 not n2870 ; n2870_not
g5013 not n2872 ; n2872_not
g5014 not n2873 ; n2873_not
g5015 not n2875 ; n2875_not
g5016 not n2876 ; n2876_not
g5017 not n2878 ; n2878_not
g5018 not n2871 ; n2871_not
g5019 not n2879 ; n2879_not
g5020 not n2881 ; n2881_not
g5021 not n2882 ; n2882_not
g5022 not n2884 ; n2884_not
g5023 not n2885 ; n2885_not
g5024 not n2887 ; n2887_not
g5025 not n2889 ; n2889_not
g5026 not n2890 ; n2890_not
g5027 not n2892 ; n2892_not
g5028 not n2893 ; n2893_not
g5029 not n2895 ; n2895_not
g5030 not n2888 ; n2888_not
g5031 not n2896 ; n2896_not
g5032 not n2898 ; n2898_not
g5033 not n2899 ; n2899_not
g5034 not n2901 ; n2901_not
g5035 not n2902 ; n2902_not
g5036 not n2904 ; n2904_not
g5037 not n2906 ; n2906_not
g5038 not n2907 ; n2907_not
g5039 not n2909 ; n2909_not
g5040 not n2910 ; n2910_not
g5041 not n2912 ; n2912_not
g5042 not n2905 ; n2905_not
g5043 not n2913 ; n2913_not
g5044 not n2915 ; n2915_not
g5045 not n2916 ; n2916_not
g5046 not n2918 ; n2918_not
g5047 not n2919 ; n2919_not
g5048 not n2921 ; n2921_not
g5049 not n2923 ; n2923_not
g5050 not n2924 ; n2924_not
g5051 not n2926 ; n2926_not
g5052 not n2927 ; n2927_not
g5053 not n2929 ; n2929_not
g5054 not n2922 ; n2922_not
g5055 not n2930 ; n2930_not
g5056 not n2932 ; n2932_not
g5057 not n2933 ; n2933_not
g5058 not n2935 ; n2935_not
g5059 not n2936 ; n2936_not
g5060 not n2938 ; n2938_not
g5061 not n2940 ; n2940_not
g5062 not n2941 ; n2941_not
g5063 not n2943 ; n2943_not
g5064 not n2944 ; n2944_not
g5065 not n2946 ; n2946_not
g5066 not n2939 ; n2939_not
g5067 not n2947 ; n2947_not
g5068 not n2949 ; n2949_not
g5069 not n2950 ; n2950_not
g5070 not n2952 ; n2952_not
g5071 not n2953 ; n2953_not
g5072 not n2955 ; n2955_not
g5073 not n2957 ; n2957_not
g5074 not n2958 ; n2958_not
g5075 not n2960 ; n2960_not
g5076 not n2961 ; n2961_not
g5077 not n2963 ; n2963_not
g5078 not n2956 ; n2956_not
g5079 not n2964 ; n2964_not
g5080 not n2966 ; n2966_not
g5081 not n2967 ; n2967_not
g5082 not n2969 ; n2969_not
g5083 not n2970 ; n2970_not
g5084 not n2972 ; n2972_not
g5085 not n2974 ; n2974_not
g5086 not n2975 ; n2975_not
g5087 not n2977 ; n2977_not
g5088 not n2978 ; n2978_not
g5089 not n2980 ; n2980_not
g5090 not n2973 ; n2973_not
g5091 not n2981 ; n2981_not
g5092 not n2983 ; n2983_not
g5093 not n2984 ; n2984_not
g5094 not n2986 ; n2986_not
g5095 not n2987 ; n2987_not
g5096 not n2989 ; n2989_not
g5097 not n2991 ; n2991_not
g5098 not n2992 ; n2992_not
g5099 not n2994 ; n2994_not
g5100 not n2995 ; n2995_not
g5101 not n2997 ; n2997_not
g5102 not n2990 ; n2990_not
g5103 not n2998 ; n2998_not
g5104 not n3000 ; n3000_not
g5105 not n3001 ; n3001_not
g5106 not n3003 ; n3003_not
g5107 not n3004 ; n3004_not
g5108 not n3006 ; n3006_not
g5109 not n3008 ; n3008_not
g5110 not n3009 ; n3009_not
g5111 not n3011 ; n3011_not
g5112 not n3012 ; n3012_not
g5113 not n3014 ; n3014_not
g5114 not n3007 ; n3007_not
g5115 not n3015 ; n3015_not
g5116 not n3017 ; n3017_not
g5117 not n3018 ; n3018_not
g5118 not n3020 ; n3020_not
g5119 not n3021 ; n3021_not
g5120 not n3023 ; n3023_not
g5121 not n3025 ; n3025_not
g5122 not n3026 ; n3026_not
g5123 not n3028 ; n3028_not
g5124 not n3029 ; n3029_not
g5125 not n3031 ; n3031_not
g5126 not n3024 ; n3024_not
g5127 not n3032 ; n3032_not
g5128 not n3034 ; n3034_not
g5129 not n3035 ; n3035_not
g5130 not n3037 ; n3037_not
g5131 not n3038 ; n3038_not
g5132 not n3040 ; n3040_not
g5133 not n3042 ; n3042_not
g5134 not n3043 ; n3043_not
g5135 not n3045 ; n3045_not
g5136 not n3046 ; n3046_not
g5137 not n3048 ; n3048_not
g5138 not n3041 ; n3041_not
g5139 not n3049 ; n3049_not
g5140 not n3051 ; n3051_not
g5141 not n3052 ; n3052_not
g5142 not n3054 ; n3054_not
g5143 not n3055 ; n3055_not
g5144 not n3057 ; n3057_not
g5145 not n3059 ; n3059_not
g5146 not n3060 ; n3060_not
g5147 not n3062 ; n3062_not
g5148 not n3063 ; n3063_not
g5149 not n3065 ; n3065_not
g5150 not n3058 ; n3058_not
g5151 not n3066 ; n3066_not
g5152 not n3068 ; n3068_not
g5153 not n3069 ; n3069_not
g5154 not n3071 ; n3071_not
g5155 not n3072 ; n3072_not
g5156 not n3074 ; n3074_not
g5157 not n3076 ; n3076_not
g5158 not n3077 ; n3077_not
g5159 not n3079 ; n3079_not
g5160 not n3080 ; n3080_not
g5161 not n3082 ; n3082_not
g5162 not n3075 ; n3075_not
g5163 not n3083 ; n3083_not
g5164 not n3085 ; n3085_not
g5165 not n3086 ; n3086_not
g5166 not n3088 ; n3088_not
g5167 not n3089 ; n3089_not
g5168 not n3091 ; n3091_not
g5169 not n3093 ; n3093_not
g5170 not n3094 ; n3094_not
g5171 not n3096 ; n3096_not
g5172 not n3097 ; n3097_not
g5173 not n3099 ; n3099_not
g5174 not n3092 ; n3092_not
g5175 not n3100 ; n3100_not
g5176 not n3102 ; n3102_not
g5177 not n3103 ; n3103_not
g5178 not n3105 ; n3105_not
g5179 not n3106 ; n3106_not
g5180 not n3108 ; n3108_not
g5181 not n3110 ; n3110_not
g5182 not n3111 ; n3111_not
g5183 not n3113 ; n3113_not
g5184 not n3114 ; n3114_not
g5185 not n3116 ; n3116_not
g5186 not n3109 ; n3109_not
g5187 not n3117 ; n3117_not
g5188 not n3119 ; n3119_not
g5189 not n3120 ; n3120_not
g5190 not n3122 ; n3122_not
g5191 not n3123 ; n3123_not
g5192 not n3125 ; n3125_not
g5193 not n3127 ; n3127_not
g5194 not n3128 ; n3128_not
g5195 not n3130 ; n3130_not
g5196 not n3131 ; n3131_not
g5197 not n3133 ; n3133_not
g5198 not n3126 ; n3126_not
g5199 not n3134 ; n3134_not
g5200 not n3136 ; n3136_not
g5201 not n3137 ; n3137_not
g5202 not n3139 ; n3139_not
g5203 not n3140 ; n3140_not
g5204 not n3142 ; n3142_not
g5205 not n3144 ; n3144_not
g5206 not n3145 ; n3145_not
g5207 not n3147 ; n3147_not
g5208 not n3148 ; n3148_not
g5209 not n3150 ; n3150_not
g5210 not n3143 ; n3143_not
g5211 not n3151 ; n3151_not
g5212 not n3153 ; n3153_not
g5213 not n3154 ; n3154_not
g5214 not n3156 ; n3156_not
g5215 not n3157 ; n3157_not
g5216 not n3159 ; n3159_not
g5217 not n3161 ; n3161_not
g5218 not n3162 ; n3162_not
g5219 not n3164 ; n3164_not
g5220 not n3165 ; n3165_not
g5221 not n3167 ; n3167_not
g5222 not n3160 ; n3160_not
g5223 not n3168 ; n3168_not
g5224 not n3170 ; n3170_not
g5225 not n3171 ; n3171_not
g5226 not n3173 ; n3173_not
g5227 not n3174 ; n3174_not
g5228 not n3176 ; n3176_not
g5229 not n3178 ; n3178_not
g5230 not n3179 ; n3179_not
g5231 not n3181 ; n3181_not
g5232 not n3182 ; n3182_not
g5233 not n3184 ; n3184_not
g5234 not n3177 ; n3177_not
g5235 not n3185 ; n3185_not
g5236 not n3187 ; n3187_not
g5237 not n3188 ; n3188_not
g5238 not n3190 ; n3190_not
g5239 not n3191 ; n3191_not
g5240 not n3193 ; n3193_not
g5241 not n3195 ; n3195_not
g5242 not n3196 ; n3196_not
g5243 not n3198 ; n3198_not
g5244 not n3199 ; n3199_not
g5245 not n3201 ; n3201_not
g5246 not n3194 ; n3194_not
g5247 not n3202 ; n3202_not
g5248 not n3204 ; n3204_not
g5249 not n3205 ; n3205_not
g5250 not n3207 ; n3207_not
g5251 not n3208 ; n3208_not
g5252 not n3210 ; n3210_not
g5253 not n3212 ; n3212_not
g5254 not n3213 ; n3213_not
g5255 not n3215 ; n3215_not
g5256 not n3216 ; n3216_not
g5257 not n3218 ; n3218_not
g5258 not n3211 ; n3211_not
g5259 not n3219 ; n3219_not
g5260 not n3221 ; n3221_not
g5261 not n3222 ; n3222_not
g5262 not n3224 ; n3224_not
g5263 not n3225 ; n3225_not
g5264 not n3227 ; n3227_not
g5265 not n3229 ; n3229_not
g5266 not n3230 ; n3230_not
g5267 not n3232 ; n3232_not
g5268 not n3233 ; n3233_not
g5269 not n3235 ; n3235_not
g5270 not n3228 ; n3228_not
g5271 not n3236 ; n3236_not
g5272 not n3238 ; n3238_not
g5273 not n3239 ; n3239_not
g5274 not n3241 ; n3241_not
g5275 not n3242 ; n3242_not
g5276 not n3244 ; n3244_not
g5277 not n3246 ; n3246_not
g5278 not n3247 ; n3247_not
g5279 not n3249 ; n3249_not
g5280 not n3250 ; n3250_not
g5281 not n3252 ; n3252_not
g5282 not n3245 ; n3245_not
g5283 not n3253 ; n3253_not
g5284 not n3255 ; n3255_not
g5285 not n3256 ; n3256_not
g5286 not n3258 ; n3258_not
g5287 not n3259 ; n3259_not
g5288 not n3261 ; n3261_not
g5289 not n3263 ; n3263_not
g5290 not n3264 ; n3264_not
g5291 not n3266 ; n3266_not
g5292 not n3267 ; n3267_not
g5293 not n3269 ; n3269_not
g5294 not n3262 ; n3262_not
g5295 not n3270 ; n3270_not
g5296 not n3272 ; n3272_not
g5297 not n3273 ; n3273_not
g5298 not n3275 ; n3275_not
g5299 not n3276 ; n3276_not
g5300 not n3278 ; n3278_not
g5301 not n3280 ; n3280_not
g5302 not n3281 ; n3281_not
g5303 not n3283 ; n3283_not
g5304 not n3284 ; n3284_not
g5305 not n3286 ; n3286_not
g5306 not n3279 ; n3279_not
g5307 not n3287 ; n3287_not
g5308 not n3289 ; n3289_not
g5309 not n3290 ; n3290_not
g5310 not n3292 ; n3292_not
g5311 not n3293 ; n3293_not
g5312 not n3295 ; n3295_not
g5313 not n3297 ; n3297_not
g5314 not n3298 ; n3298_not
g5315 not n3300 ; n3300_not
g5316 not n3301 ; n3301_not
g5317 not n3303 ; n3303_not
g5318 not n3296 ; n3296_not
g5319 not n3304 ; n3304_not
g5320 not n3306 ; n3306_not
g5321 not n3307 ; n3307_not
g5322 not n3309 ; n3309_not
g5323 not n3310 ; n3310_not
g5324 not n3312 ; n3312_not
g5325 not n3314 ; n3314_not
g5326 not n3315 ; n3315_not
g5327 not n3317 ; n3317_not
g5328 not n3318 ; n3318_not
g5329 not n3320 ; n3320_not
g5330 not n3313 ; n3313_not
g5331 not n3321 ; n3321_not
g5332 not n3323 ; n3323_not
g5333 not n3324 ; n3324_not
g5334 not n3326 ; n3326_not
g5335 not n3327 ; n3327_not
g5336 not n3329 ; n3329_not
g5337 not n3331 ; n3331_not
g5338 not n3332 ; n3332_not
g5339 not n3334 ; n3334_not
g5340 not n3335 ; n3335_not
g5341 not n3337 ; n3337_not
g5342 not n3330 ; n3330_not
g5343 not n3338 ; n3338_not
g5344 not n3340 ; n3340_not
g5345 not n3341 ; n3341_not
g5346 not n3343 ; n3343_not
g5347 not n3344 ; n3344_not
g5348 not n3346 ; n3346_not
g5349 not n3348 ; n3348_not
g5350 not n3349 ; n3349_not
g5351 not n3351 ; n3351_not
g5352 not n3352 ; n3352_not
g5353 not n3354 ; n3354_not
g5354 not n3347 ; n3347_not
g5355 not n3355 ; n3355_not
g5356 not n3357 ; n3357_not
g5357 not n3358 ; n3358_not
g5358 not n3360 ; n3360_not
g5359 not n3361 ; n3361_not
g5360 not n3363 ; n3363_not
g5361 not n3365 ; n3365_not
g5362 not n3366 ; n3366_not
g5363 not n3368 ; n3368_not
g5364 not n3369 ; n3369_not
g5365 not n3371 ; n3371_not
g5366 not n3364 ; n3364_not
g5367 not n3372 ; n3372_not
g5368 not n3374 ; n3374_not
g5369 not n3375 ; n3375_not
g5370 not n3377 ; n3377_not
g5371 not n3378 ; n3378_not
g5372 not n3380 ; n3380_not
g5373 not n3382 ; n3382_not
g5374 not n3383 ; n3383_not
g5375 not n3385 ; n3385_not
g5376 not n3386 ; n3386_not
g5377 not n3388 ; n3388_not
g5378 not n3381 ; n3381_not
g5379 not n3389 ; n3389_not
g5380 not n3391 ; n3391_not
g5381 not n3392 ; n3392_not
g5382 not n3394 ; n3394_not
g5383 not n3395 ; n3395_not
g5384 not n3397 ; n3397_not
g5385 not n3399 ; n3399_not
g5386 not n3400 ; n3400_not
g5387 not n3402 ; n3402_not
g5388 not n3403 ; n3403_not
g5389 not n3405 ; n3405_not
g5390 not n3398 ; n3398_not
g5391 not n3406 ; n3406_not
g5392 not n3408 ; n3408_not
g5393 not n3409 ; n3409_not
g5394 not n3411 ; n3411_not
g5395 not n3412 ; n3412_not
g5396 not n3414 ; n3414_not
g5397 not n3415 ; n3415_not
g5398 not n3417 ; n3417_not
g5399 not n3418 ; n3418_not
g5400 not n3420 ; n3420_not
g5401 not n3421 ; n3421_not
g5402 not n3423 ; n3423_not
g5403 not n3424 ; n3424_not
g5404 not n3426 ; n3426_not
g5405 not n3427 ; n3427_not
g5406 not n3429 ; n3429_not
g5407 not n3430 ; n3430_not
g5408 not n3432 ; n3432_not
g5409 not n3433 ; n3433_not
g5410 not n3435 ; n3435_not
g5411 not n3436 ; n3436_not
g5412 not n3438 ; n3438_not
g5413 not n3439 ; n3439_not
g5414 not n3441 ; n3441_not
g5415 not n3442 ; n3442_not
g5416 not n3444 ; n3444_not
g5417 not n3445 ; n3445_not
g5418 not n3447 ; n3447_not
g5419 not n3448 ; n3448_not
g5420 not n3450 ; n3450_not
g5421 not n3451 ; n3451_not
g5422 not n3453 ; n3453_not
g5423 not n3454 ; n3454_not
g5424 not n3456 ; n3456_not
g5425 not n3457 ; n3457_not
g5426 not n3459 ; n3459_not
g5427 not n3460 ; n3460_not
g5428 not n3462 ; n3462_not
g5429 not n3463 ; n3463_not
g5430 not n3465 ; n3465_not
g5431 not n3466 ; n3466_not
g5432 not n3468 ; n3468_not
g5433 not n3469 ; n3469_not
g5434 not n3471 ; n3471_not
g5435 not n3472 ; n3472_not
g5436 not n3474 ; n3474_not
g5437 not n3475 ; n3475_not
g5438 not n3477 ; n3477_not
g5439 not n3478 ; n3478_not
g5440 not n3480 ; n3480_not
g5441 not n3481 ; n3481_not
g5442 not n3483 ; n3483_not
g5443 not n3484 ; n3484_not
g5444 not n3486 ; n3486_not
g5445 not n3487 ; n3487_not
g5446 not n3489 ; n3489_not
g5447 not n3490 ; n3490_not
g5448 not n3492 ; n3492_not
g5449 not n3493 ; n3493_not
g5450 not n3495 ; n3495_not
g5451 not n3496 ; n3496_not
g5452 not n3498 ; n3498_not
g5453 not n3499 ; n3499_not
g5454 not n3501 ; n3501_not
g5455 not n3502 ; n3502_not
g5456 not n3504 ; n3504_not
g5457 not n3505 ; n3505_not
g5458 not n3507 ; n3507_not
g5459 not n3508 ; n3508_not
g5460 not n3510 ; n3510_not
g5461 not n3511 ; n3511_not
g5462 not n3513 ; n3513_not
g5463 not n3514 ; n3514_not
g5464 not n3516 ; n3516_not
g5465 not n3517 ; n3517_not
g5466 not n3519 ; n3519_not
g5467 not n3520 ; n3520_not
g5468 not n3522 ; n3522_not
g5469 not n3523 ; n3523_not
g5470 not n3525 ; n3525_not
g5471 not n3526 ; n3526_not
g5472 not n3528 ; n3528_not
g5473 not n3529 ; n3529_not
g5474 not n3531 ; n3531_not
g5475 not n3532 ; n3532_not
g5476 not n3534 ; n3534_not
g5477 not n3535 ; n3535_not
g5478 not n3537 ; n3537_not
g5479 not n3538 ; n3538_not
g5480 not n3540 ; n3540_not
g5481 not n3541 ; n3541_not
g5482 not n3543 ; n3543_not
g5483 not n3544 ; n3544_not
g5484 not n3546 ; n3546_not
g5485 not n3547 ; n3547_not
g5486 not n3549 ; n3549_not
g5487 not n3550 ; n3550_not
g5488 not n3552 ; n3552_not
g5489 not n3553 ; n3553_not
g5490 not n3555 ; n3555_not
g5491 not n3556 ; n3556_not
g5492 not n3558 ; n3558_not
g5493 not n3559 ; n3559_not
g5494 not n3561 ; n3561_not
g5495 not n3562 ; n3562_not
g5496 not n3564 ; n3564_not
g5497 not n3565 ; n3565_not
g5498 not n3567 ; n3567_not
g5499 not n3568 ; n3568_not
g5500 not n3570 ; n3570_not
g5501 not n3571 ; n3571_not
g5502 not n3573 ; n3573_not
g5503 not n3574 ; n3574_not
g5504 not n3576 ; n3576_not
g5505 not n3577 ; n3577_not
g5506 not n3579 ; n3579_not
g5507 not n3580 ; n3580_not
g5508 not n3582 ; n3582_not
g5509 not n3583 ; n3583_not
g5510 not n3585 ; n3585_not
g5511 not n3586 ; n3586_not
g5512 not n3588 ; n3588_not
g5513 not n3589 ; n3589_not
g5514 not n3591 ; n3591_not
g5515 not n3592 ; n3592_not
g5516 not n3594 ; n3594_not
g5517 not n3595 ; n3595_not
g5518 not n3597 ; n3597_not
g5519 not n3598 ; n3598_not
o result[0]
o result[1]
o result[2]
o result[3]
o result[4]
o result[5]
o result[6]
o result[7]
o result[8]
o result[9]
o result[10]
o result[11]
o result[12]
o result[13]
o result[14]
o result[15]
o result[16]
o result[17]
o result[18]
o result[19]
o result[20]
o result[21]
o result[22]
o result[23]
o result[24]
o result[25]
o result[26]
o result[27]
o result[28]
o result[29]
o result[30]
o result[31]
o result[32]
o result[33]
o result[34]
o result[35]
o result[36]
o result[37]
o result[38]
o result[39]
o result[40]
o result[41]
o result[42]
o result[43]
o result[44]
o result[45]
o result[46]
o result[47]
o result[48]
o result[49]
o result[50]
o result[51]
o result[52]
o result[53]
o result[54]
o result[55]
o result[56]
o result[57]
o result[58]
o result[59]
o result[60]
o result[61]
o result[62]
o result[63]
o result[64]
o result[65]
o result[66]
o result[67]
o result[68]
o result[69]
o result[70]
o result[71]
o result[72]
o result[73]
o result[74]
o result[75]
o result[76]
o result[77]
o result[78]
o result[79]
o result[80]
o result[81]
o result[82]
o result[83]
o result[84]
o result[85]
o result[86]
o result[87]
o result[88]
o result[89]
o result[90]
o result[91]
o result[92]
o result[93]
o result[94]
o result[95]
o result[96]
o result[97]
o result[98]
o result[99]
o result[100]
o result[101]
o result[102]
o result[103]
o result[104]
o result[105]
o result[106]
o result[107]
o result[108]
o result[109]
o result[110]
o result[111]
o result[112]
o result[113]
o result[114]
o result[115]
o result[116]
o result[117]
o result[118]
o result[119]
o result[120]
o result[121]
o result[122]
o result[123]
o result[124]
o result[125]
o result[126]
o result[127]
