name max
i in0[0]
i in0[1]
i in0[2]
i in0[3]
i in0[4]
i in0[5]
i in0[6]
i in0[7]
i in0[8]
i in0[9]
i in0[10]
i in0[11]
i in0[12]
i in0[13]
i in0[14]
i in0[15]
i in0[16]
i in0[17]
i in0[18]
i in0[19]
i in0[20]
i in0[21]
i in0[22]
i in0[23]
i in0[24]
i in0[25]
i in0[26]
i in0[27]
i in0[28]
i in0[29]
i in0[30]
i in0[31]
i in0[32]
i in0[33]
i in0[34]
i in0[35]
i in0[36]
i in0[37]
i in0[38]
i in0[39]
i in0[40]
i in0[41]
i in0[42]
i in0[43]
i in0[44]
i in0[45]
i in0[46]
i in0[47]
i in0[48]
i in0[49]
i in0[50]
i in0[51]
i in0[52]
i in0[53]
i in0[54]
i in0[55]
i in0[56]
i in0[57]
i in0[58]
i in0[59]
i in0[60]
i in0[61]
i in0[62]
i in0[63]
i in0[64]
i in0[65]
i in0[66]
i in0[67]
i in0[68]
i in0[69]
i in0[70]
i in0[71]
i in0[72]
i in0[73]
i in0[74]
i in0[75]
i in0[76]
i in0[77]
i in0[78]
i in0[79]
i in0[80]
i in0[81]
i in0[82]
i in0[83]
i in0[84]
i in0[85]
i in0[86]
i in0[87]
i in0[88]
i in0[89]
i in0[90]
i in0[91]
i in0[92]
i in0[93]
i in0[94]
i in0[95]
i in0[96]
i in0[97]
i in0[98]
i in0[99]
i in0[100]
i in0[101]
i in0[102]
i in0[103]
i in0[104]
i in0[105]
i in0[106]
i in0[107]
i in0[108]
i in0[109]
i in0[110]
i in0[111]
i in0[112]
i in0[113]
i in0[114]
i in0[115]
i in0[116]
i in0[117]
i in0[118]
i in0[119]
i in0[120]
i in0[121]
i in0[122]
i in0[123]
i in0[124]
i in0[125]
i in0[126]
i in0[127]
i in1[0]
i in1[1]
i in1[2]
i in1[3]
i in1[4]
i in1[5]
i in1[6]
i in1[7]
i in1[8]
i in1[9]
i in1[10]
i in1[11]
i in1[12]
i in1[13]
i in1[14]
i in1[15]
i in1[16]
i in1[17]
i in1[18]
i in1[19]
i in1[20]
i in1[21]
i in1[22]
i in1[23]
i in1[24]
i in1[25]
i in1[26]
i in1[27]
i in1[28]
i in1[29]
i in1[30]
i in1[31]
i in1[32]
i in1[33]
i in1[34]
i in1[35]
i in1[36]
i in1[37]
i in1[38]
i in1[39]
i in1[40]
i in1[41]
i in1[42]
i in1[43]
i in1[44]
i in1[45]
i in1[46]
i in1[47]
i in1[48]
i in1[49]
i in1[50]
i in1[51]
i in1[52]
i in1[53]
i in1[54]
i in1[55]
i in1[56]
i in1[57]
i in1[58]
i in1[59]
i in1[60]
i in1[61]
i in1[62]
i in1[63]
i in1[64]
i in1[65]
i in1[66]
i in1[67]
i in1[68]
i in1[69]
i in1[70]
i in1[71]
i in1[72]
i in1[73]
i in1[74]
i in1[75]
i in1[76]
i in1[77]
i in1[78]
i in1[79]
i in1[80]
i in1[81]
i in1[82]
i in1[83]
i in1[84]
i in1[85]
i in1[86]
i in1[87]
i in1[88]
i in1[89]
i in1[90]
i in1[91]
i in1[92]
i in1[93]
i in1[94]
i in1[95]
i in1[96]
i in1[97]
i in1[98]
i in1[99]
i in1[100]
i in1[101]
i in1[102]
i in1[103]
i in1[104]
i in1[105]
i in1[106]
i in1[107]
i in1[108]
i in1[109]
i in1[110]
i in1[111]
i in1[112]
i in1[113]
i in1[114]
i in1[115]
i in1[116]
i in1[117]
i in1[118]
i in1[119]
i in1[120]
i in1[121]
i in1[122]
i in1[123]
i in1[124]
i in1[125]
i in1[126]
i in1[127]
i in2[0]
i in2[1]
i in2[2]
i in2[3]
i in2[4]
i in2[5]
i in2[6]
i in2[7]
i in2[8]
i in2[9]
i in2[10]
i in2[11]
i in2[12]
i in2[13]
i in2[14]
i in2[15]
i in2[16]
i in2[17]
i in2[18]
i in2[19]
i in2[20]
i in2[21]
i in2[22]
i in2[23]
i in2[24]
i in2[25]
i in2[26]
i in2[27]
i in2[28]
i in2[29]
i in2[30]
i in2[31]
i in2[32]
i in2[33]
i in2[34]
i in2[35]
i in2[36]
i in2[37]
i in2[38]
i in2[39]
i in2[40]
i in2[41]
i in2[42]
i in2[43]
i in2[44]
i in2[45]
i in2[46]
i in2[47]
i in2[48]
i in2[49]
i in2[50]
i in2[51]
i in2[52]
i in2[53]
i in2[54]
i in2[55]
i in2[56]
i in2[57]
i in2[58]
i in2[59]
i in2[60]
i in2[61]
i in2[62]
i in2[63]
i in2[64]
i in2[65]
i in2[66]
i in2[67]
i in2[68]
i in2[69]
i in2[70]
i in2[71]
i in2[72]
i in2[73]
i in2[74]
i in2[75]
i in2[76]
i in2[77]
i in2[78]
i in2[79]
i in2[80]
i in2[81]
i in2[82]
i in2[83]
i in2[84]
i in2[85]
i in2[86]
i in2[87]
i in2[88]
i in2[89]
i in2[90]
i in2[91]
i in2[92]
i in2[93]
i in2[94]
i in2[95]
i in2[96]
i in2[97]
i in2[98]
i in2[99]
i in2[100]
i in2[101]
i in2[102]
i in2[103]
i in2[104]
i in2[105]
i in2[106]
i in2[107]
i in2[108]
i in2[109]
i in2[110]
i in2[111]
i in2[112]
i in2[113]
i in2[114]
i in2[115]
i in2[116]
i in2[117]
i in2[118]
i in2[119]
i in2[120]
i in2[121]
i in2[122]
i in2[123]
i in2[124]
i in2[125]
i in2[126]
i in2[127]
i in3[0]
i in3[1]
i in3[2]
i in3[3]
i in3[4]
i in3[5]
i in3[6]
i in3[7]
i in3[8]
i in3[9]
i in3[10]
i in3[11]
i in3[12]
i in3[13]
i in3[14]
i in3[15]
i in3[16]
i in3[17]
i in3[18]
i in3[19]
i in3[20]
i in3[21]
i in3[22]
i in3[23]
i in3[24]
i in3[25]
i in3[26]
i in3[27]
i in3[28]
i in3[29]
i in3[30]
i in3[31]
i in3[32]
i in3[33]
i in3[34]
i in3[35]
i in3[36]
i in3[37]
i in3[38]
i in3[39]
i in3[40]
i in3[41]
i in3[42]
i in3[43]
i in3[44]
i in3[45]
i in3[46]
i in3[47]
i in3[48]
i in3[49]
i in3[50]
i in3[51]
i in3[52]
i in3[53]
i in3[54]
i in3[55]
i in3[56]
i in3[57]
i in3[58]
i in3[59]
i in3[60]
i in3[61]
i in3[62]
i in3[63]
i in3[64]
i in3[65]
i in3[66]
i in3[67]
i in3[68]
i in3[69]
i in3[70]
i in3[71]
i in3[72]
i in3[73]
i in3[74]
i in3[75]
i in3[76]
i in3[77]
i in3[78]
i in3[79]
i in3[80]
i in3[81]
i in3[82]
i in3[83]
i in3[84]
i in3[85]
i in3[86]
i in3[87]
i in3[88]
i in3[89]
i in3[90]
i in3[91]
i in3[92]
i in3[93]
i in3[94]
i in3[95]
i in3[96]
i in3[97]
i in3[98]
i in3[99]
i in3[100]
i in3[101]
i in3[102]
i in3[103]
i in3[104]
i in3[105]
i in3[106]
i in3[107]
i in3[108]
i in3[109]
i in3[110]
i in3[111]
i in3[112]
i in3[113]
i in3[114]
i in3[115]
i in3[116]
i in3[117]
i in3[118]
i in3[119]
i in3[120]
i in3[121]
i in3[122]
i in3[123]
i in3[124]
i in3[125]
i in3[126]
i in3[127]

g1 and in2[119] in3[119]_not ; n643
g2 and in2[119]_not in3[119] ; n644
g3 and in2[118]_not in3[118] ; n645
g4 and n644_not n645_not ; n646
g5 and in2[117]_not in3[117] ; n647
g6 and in2[116] in3[116]_not ; n648
g7 and n647_not n648 ; n649
g8 and in2[117] in3[117]_not ; n650
g9 and n649_not n650_not ; n651
g10 and n646 n651_not ; n652
g11 and in3[118]_not n644_not ; n653
g12 and in2[118] n653 ; n654
g13 and in2[112]_not in3[112] ; n655
g14 and in2[115]_not in3[115] ; n656
g15 and in2[114]_not in3[114] ; n657
g16 and n656_not n657_not ; n658
g17 and in2[113]_not in3[113] ; n659
g18 and in2[111] in3[111]_not ; n660
g19 and in2[111]_not in3[111] ; n661
g20 and in2[110]_not in3[110] ; n662
g21 and n661_not n662_not ; n663
g22 and in2[109]_not in3[109] ; n664
g23 and in2[108] in3[108]_not ; n665
g24 and n664_not n665 ; n666
g25 and in2[109] in3[109]_not ; n667
g26 and n666_not n667_not ; n668
g27 and n663 n668_not ; n669
g28 and in3[110]_not n661_not ; n670
g29 and in2[110] n670 ; n671
g30 and in2[103] in3[103]_not ; n672
g31 and in2[103]_not in3[103] ; n673
g32 and in2[102]_not in3[102] ; n674
g33 and n673_not n674_not ; n675
g34 and in2[101]_not in3[101] ; n676
g35 and in2[100] in3[100]_not ; n677
g36 and n676_not n677 ; n678
g37 and in2[101] in3[101]_not ; n679
g38 and n678_not n679_not ; n680
g39 and n675 n680_not ; n681
g40 and in3[102]_not n673_not ; n682
g41 and in2[102] n682 ; n683
g42 and in2[96]_not in3[96] ; n684
g43 and in2[99]_not in3[99] ; n685
g44 and in2[98]_not in3[98] ; n686
g45 and n685_not n686_not ; n687
g46 and in2[97]_not in3[97] ; n688
g47 and in2[95] in3[95]_not ; n689
g48 and in2[95]_not in3[95] ; n690
g49 and in2[94]_not in3[94] ; n691
g50 and n690_not n691_not ; n692
g51 and in2[93]_not in3[93] ; n693
g52 and in2[92] in3[92]_not ; n694
g53 and n693_not n694 ; n695
g54 and in2[93] in3[93]_not ; n696
g55 and n695_not n696_not ; n697
g56 and n692 n697_not ; n698
g57 and in3[94]_not n690_not ; n699
g58 and in2[94] n699 ; n700
g59 and in2[87] in3[87]_not ; n701
g60 and in2[87]_not in3[87] ; n702
g61 and in2[86]_not in3[86] ; n703
g62 and n702_not n703_not ; n704
g63 and in2[85]_not in3[85] ; n705
g64 and in2[84] in3[84]_not ; n706
g65 and n705_not n706 ; n707
g66 and in2[85] in3[85]_not ; n708
g67 and n707_not n708_not ; n709
g68 and n704 n709_not ; n710
g69 and in3[86]_not n702_not ; n711
g70 and in2[86] n711 ; n712
g71 and in2[80]_not in3[80] ; n713
g72 and in2[83]_not in3[83] ; n714
g73 and in2[82]_not in3[82] ; n715
g74 and n714_not n715_not ; n716
g75 and in2[81]_not in3[81] ; n717
g76 and in2[79] in3[79]_not ; n718
g77 and in2[79]_not in3[79] ; n719
g78 and in2[78]_not in3[78] ; n720
g79 and n719_not n720_not ; n721
g80 and in2[77]_not in3[77] ; n722
g81 and in2[76] in3[76]_not ; n723
g82 and n722_not n723 ; n724
g83 and in2[77] in3[77]_not ; n725
g84 and n724_not n725_not ; n726
g85 and n721 n726_not ; n727
g86 and in3[78]_not n719_not ; n728
g87 and in2[78] n728 ; n729
g88 and in2[71] in3[71]_not ; n730
g89 and in2[71]_not in3[71] ; n731
g90 and in2[70]_not in3[70] ; n732
g91 and n731_not n732_not ; n733
g92 and in2[69]_not in3[69] ; n734
g93 and in2[68] in3[68]_not ; n735
g94 and n734_not n735 ; n736
g95 and in2[69] in3[69]_not ; n737
g96 and n736_not n737_not ; n738
g97 and n733 n738_not ; n739
g98 and in3[70]_not n731_not ; n740
g99 and in2[70] n740 ; n741
g100 and in2[67]_not in3[67] ; n742
g101 and in2[66]_not in3[66] ; n743
g102 and n742_not n743_not ; n744
g103 and in2[65]_not in3[65] ; n745
g104 and in2[63] in3[63]_not ; n746
g105 and in2[63]_not in3[63] ; n747
g106 and in2[62]_not in3[62] ; n748
g107 and n747_not n748_not ; n749
g108 and in2[60]_not in3[60] ; n750
g109 and in2[61]_not in3[61] ; n751
g110 and n750_not n751_not ; n752
g111 and n749 n752 ; n753
g112 and in2[59] in3[59]_not ; n754
g113 and in2[59]_not in3[59] ; n755
g114 and in2[58]_not in3[58] ; n756
g115 and n755_not n756_not ; n757
g116 and in2[57]_not in3[57] ; n758
g117 and in2[56] in3[56]_not ; n759
g118 and n758_not n759 ; n760
g119 and in2[57] in3[57]_not ; n761
g120 and n760_not n761_not ; n762
g121 and in2[58] in3[58]_not ; n763
g122 and n762 n763_not ; n764
g123 and n757 n764_not ; n765
g124 and n754_not n765_not ; n766
g125 and n753 n766_not ; n767
g126 and in2[60] in3[60]_not ; n768
g127 and n751_not n768 ; n769
g128 and in2[61] in3[61]_not ; n770
g129 and n769_not n770_not ; n771
g130 and n749 n771_not ; n772
g131 and in3[62]_not n747_not ; n773
g132 and in2[62] n773 ; n774
g133 and in2[47] in3[47]_not ; n775
g134 and in2[47]_not in3[47] ; n776
g135 and in2[46]_not in3[46] ; n777
g136 and n776_not n777_not ; n778
g137 and in2[44]_not in3[44] ; n779
g138 and in2[45]_not in3[45] ; n780
g139 and n779_not n780_not ; n781
g140 and n778 n781 ; n782
g141 and in2[43] in3[43]_not ; n783
g142 and in2[43]_not in3[43] ; n784
g143 and in2[42]_not in3[42] ; n785
g144 and n784_not n785_not ; n786
g145 and in2[41]_not in3[41] ; n787
g146 and in2[40] in3[40]_not ; n788
g147 and n787_not n788 ; n789
g148 and in2[41] in3[41]_not ; n790
g149 and n789_not n790_not ; n791
g150 and in2[42] in3[42]_not ; n792
g151 and n791 n792_not ; n793
g152 and n786 n793_not ; n794
g153 and n783_not n794_not ; n795
g154 and n782 n795_not ; n796
g155 and in2[44] in3[44]_not ; n797
g156 and n780_not n797 ; n798
g157 and in2[45] in3[45]_not ; n799
g158 and n798_not n799_not ; n800
g159 and n778 n800_not ; n801
g160 and in3[46]_not n776_not ; n802
g161 and in2[46] n802 ; n803
g162 and in2[32]_not in3[32] ; n804
g163 and in2[31]_not in3[31] ; n805
g164 and in2[30]_not in3[30] ; n806
g165 and in2[29]_not in3[29] ; n807
g166 and in2[28]_not in3[28] ; n808
g167 and in2[27]_not in3[27] ; n809
g168 and in2[26]_not in3[26] ; n810
g169 and in2[23]_not in3[23] ; n811
g170 and in2[22]_not in3[22] ; n812
g171 and in2[21]_not in3[21] ; n813
g172 and in2[20]_not in3[20] ; n814
g173 and in2[19]_not in3[19] ; n815
g174 and in2[18]_not in3[18] ; n816
g175 and in2[15]_not in3[15] ; n817
g176 and in2[14]_not in3[14] ; n818
g177 and in2[13]_not in3[13] ; n819
g178 and in2[12]_not in3[12] ; n820
g179 and in2[11]_not in3[11] ; n821
g180 and in2[10]_not in3[10] ; n822
g181 and in2[7]_not in3[7] ; n823
g182 and in2[6]_not in3[6] ; n824
g183 and in2[3]_not in3[3] ; n825
g184 and in2[0] in3[0]_not ; n826
g185 and in2[1] n826 ; n827
g186 and in3[1] n827_not ; n828
g187 and in2[2]_not in3[2] ; n829
g188 and in2[1]_not n826_not ; n830
g189 and n829_not n830_not ; n831
g190 and n828_not n831 ; n832
g191 and in2[2] in3[2]_not ; n833
g192 and n832_not n833_not ; n834
g193 and n825_not n834_not ; n835
g194 and in2[3] in3[3]_not ; n836
g195 and n835_not n836_not ; n837
g196 and in2[4]_not n837 ; n838
g197 and in3[4]_not n838_not ; n839
g198 and in2[4] n837_not ; n840
g199 and n839_not n840_not ; n841
g200 and in2[5]_not n841 ; n842
g201 and in3[5]_not n842_not ; n843
g202 and in2[5] n841_not ; n844
g203 and n843_not n844_not ; n845
g204 and n824_not n845_not ; n846
g205 and in2[6] in3[6]_not ; n847
g206 and n846_not n847_not ; n848
g207 and n823_not n848_not ; n849
g208 and in2[7] in3[7]_not ; n850
g209 and n849_not n850_not ; n851
g210 and in2[8]_not n851 ; n852
g211 and in3[8]_not n852_not ; n853
g212 and in2[8] n851_not ; n854
g213 and n853_not n854_not ; n855
g214 and in2[9]_not n855 ; n856
g215 and in3[9]_not n856_not ; n857
g216 and in2[9] n855_not ; n858
g217 and n857_not n858_not ; n859
g218 and n822_not n859_not ; n860
g219 and in2[10] in3[10]_not ; n861
g220 and n860_not n861_not ; n862
g221 and n821_not n862_not ; n863
g222 and in2[11] in3[11]_not ; n864
g223 and n863_not n864_not ; n865
g224 and n820_not n865_not ; n866
g225 and in2[12] in3[12]_not ; n867
g226 and n866_not n867_not ; n868
g227 and n819_not n868_not ; n869
g228 and in2[13] in3[13]_not ; n870
g229 and n869_not n870_not ; n871
g230 and n818_not n871_not ; n872
g231 and in2[14] in3[14]_not ; n873
g232 and n872_not n873_not ; n874
g233 and n817_not n874_not ; n875
g234 and in2[15] in3[15]_not ; n876
g235 and n875_not n876_not ; n877
g236 and in2[16]_not n877 ; n878
g237 and in3[16]_not n878_not ; n879
g238 and in2[16] n877_not ; n880
g239 and n879_not n880_not ; n881
g240 and in2[17]_not n881 ; n882
g241 and in3[17]_not n882_not ; n883
g242 and in2[17] n881_not ; n884
g243 and n883_not n884_not ; n885
g244 and n816_not n885_not ; n886
g245 and in2[18] in3[18]_not ; n887
g246 and n886_not n887_not ; n888
g247 and n815_not n888_not ; n889
g248 and in2[19] in3[19]_not ; n890
g249 and n889_not n890_not ; n891
g250 and n814_not n891_not ; n892
g251 and in2[20] in3[20]_not ; n893
g252 and n892_not n893_not ; n894
g253 and n813_not n894_not ; n895
g254 and in2[21] in3[21]_not ; n896
g255 and n895_not n896_not ; n897
g256 and n812_not n897_not ; n898
g257 and in2[22] in3[22]_not ; n899
g258 and n898_not n899_not ; n900
g259 and n811_not n900_not ; n901
g260 and in2[23] in3[23]_not ; n902
g261 and n901_not n902_not ; n903
g262 and in2[24]_not n903 ; n904
g263 and in3[24]_not n904_not ; n905
g264 and in2[24] n903_not ; n906
g265 and n905_not n906_not ; n907
g266 and in2[25]_not n907 ; n908
g267 and in3[25]_not n908_not ; n909
g268 and in2[25] n907_not ; n910
g269 and n909_not n910_not ; n911
g270 and n810_not n911_not ; n912
g271 and in2[26] in3[26]_not ; n913
g272 and n912_not n913_not ; n914
g273 and n809_not n914_not ; n915
g274 and in2[27] in3[27]_not ; n916
g275 and n915_not n916_not ; n917
g276 and n808_not n917_not ; n918
g277 and in2[28] in3[28]_not ; n919
g278 and n918_not n919_not ; n920
g279 and n807_not n920_not ; n921
g280 and in2[29] in3[29]_not ; n922
g281 and n921_not n922_not ; n923
g282 and n806_not n923_not ; n924
g283 and in2[30] in3[30]_not ; n925
g284 and n924_not n925_not ; n926
g285 and n805_not n926_not ; n927
g286 and in2[31] in3[31]_not ; n928
g287 and n927_not n928_not ; n929
g288 and in2[39]_not in3[39] ; n930
g289 and in2[38]_not in3[38] ; n931
g290 and n930_not n931_not ; n932
g291 and in2[36]_not in3[36] ; n933
g292 and in2[37]_not in3[37] ; n934
g293 and n933_not n934_not ; n935
g294 and n932 n935 ; n936
g295 and in2[33]_not in3[33] ; n937
g296 and in2[35]_not in3[35] ; n938
g297 and in2[34]_not in3[34] ; n939
g298 and n938_not n939_not ; n940
g299 and n937_not n940 ; n941
g300 and n936 n941 ; n942
g301 and n929_not n942 ; n943
g302 and n804_not n943 ; n944
g303 and in2[39] in3[39]_not ; n945
g304 and in2[36] in3[36]_not ; n946
g305 and n934_not n946 ; n947
g306 and in2[37] in3[37]_not ; n948
g307 and n947_not n948_not ; n949
g308 and n932 n949_not ; n950
g309 and in3[38]_not n930_not ; n951
g310 and in2[38] n951 ; n952
g311 and in2[35] in3[35]_not ; n953
g312 and in3[32]_not n937_not ; n954
g313 and in2[32] n954 ; n955
g314 and in2[33] in3[33]_not ; n956
g315 and n955_not n956_not ; n957
g316 and in2[34] in3[34]_not ; n958
g317 and n957 n958_not ; n959
g318 and n940 n959_not ; n960
g319 and n953_not n960_not ; n961
g320 and n936 n961_not ; n962
g321 and n952_not n962_not ; n963
g322 and n950_not n963 ; n964
g323 and n945_not n964 ; n965
g324 and n944_not n965 ; n966
g325 and in2[40]_not in3[40] ; n967
g326 and n787_not n967_not ; n968
g327 and n786 n968 ; n969
g328 and n782 n969 ; n970
g329 and n966_not n970 ; n971
g330 and n803_not n971_not ; n972
g331 and n801_not n972 ; n973
g332 and n796_not n973 ; n974
g333 and n775_not n974 ; n975
g334 and in2[48]_not in3[48] ; n976
g335 and in2[55]_not in3[55] ; n977
g336 and in2[54]_not in3[54] ; n978
g337 and n977_not n978_not ; n979
g338 and in2[53]_not in3[53] ; n980
g339 and in2[52]_not in3[52] ; n981
g340 and n980_not n981_not ; n982
g341 and n979 n982 ; n983
g342 and in2[49]_not in3[49] ; n984
g343 and in2[51]_not in3[51] ; n985
g344 and in2[50]_not in3[50] ; n986
g345 and n985_not n986_not ; n987
g346 and n984_not n987 ; n988
g347 and n983 n988 ; n989
g348 and n976_not n989 ; n990
g349 and n975_not n990 ; n991
g350 and in2[55] in3[55]_not ; n992
g351 and in2[51] in3[51]_not ; n993
g352 and in3[48]_not n984_not ; n994
g353 and in2[48] n994 ; n995
g354 and in2[49] in3[49]_not ; n996
g355 and n995_not n996_not ; n997
g356 and in2[50] in3[50]_not ; n998
g357 and n997 n998_not ; n999
g358 and n987 n999_not ; n1000
g359 and n993_not n1000_not ; n1001
g360 and n983 n1001_not ; n1002
g361 and in2[52] in3[52]_not ; n1003
g362 and n980_not n1003 ; n1004
g363 and in2[53] in3[53]_not ; n1005
g364 and n1004_not n1005_not ; n1006
g365 and in2[54] in3[54]_not ; n1007
g366 and n1006 n1007_not ; n1008
g367 and n979 n1008_not ; n1009
g368 and n1002_not n1009_not ; n1010
g369 and n992_not n1010 ; n1011
g370 and n991_not n1011 ; n1012
g371 and in2[56]_not in3[56] ; n1013
g372 and n758_not n1013_not ; n1014
g373 and n753 n1014 ; n1015
g374 and n757 n1015 ; n1016
g375 and n1012_not n1016 ; n1017
g376 and n774_not n1017_not ; n1018
g377 and n772_not n1018 ; n1019
g378 and n767_not n1019 ; n1020
g379 and n746_not n1020 ; n1021
g380 and in2[64]_not in3[64] ; n1022
g381 and n1021_not n1022_not ; n1023
g382 and n745_not n1023 ; n1024
g383 and n744 n1024 ; n1025
g384 and in2[67] in3[67]_not ; n1026
g385 and in2[64] in3[64]_not ; n1027
g386 and n745_not n1027 ; n1028
g387 and in2[65] in3[65]_not ; n1029
g388 and n1028_not n1029_not ; n1030
g389 and in2[66] in3[66]_not ; n1031
g390 and n1030 n1031_not ; n1032
g391 and n744 n1032_not ; n1033
g392 and n1026_not n1033_not ; n1034
g393 and n1025_not n1034 ; n1035
g394 and in2[68]_not in3[68] ; n1036
g395 and n734_not n1036_not ; n1037
g396 and n733 n1037 ; n1038
g397 and n1035_not n1038 ; n1039
g398 and n741_not n1039_not ; n1040
g399 and n739_not n1040 ; n1041
g400 and n730_not n1041 ; n1042
g401 and in2[75]_not in3[75] ; n1043
g402 and in2[74]_not in3[74] ; n1044
g403 and n1043_not n1044_not ; n1045
g404 and in2[73]_not in3[73] ; n1046
g405 and in2[72]_not in3[72] ; n1047
g406 and n1046_not n1047_not ; n1048
g407 and n1045 n1048 ; n1049
g408 and n1042_not n1049 ; n1050
g409 and in2[75] in3[75]_not ; n1051
g410 and in2[72] in3[72]_not ; n1052
g411 and n1046_not n1052 ; n1053
g412 and in2[73] in3[73]_not ; n1054
g413 and n1053_not n1054_not ; n1055
g414 and in2[74] in3[74]_not ; n1056
g415 and n1055 n1056_not ; n1057
g416 and n1045 n1057_not ; n1058
g417 and n1051_not n1058_not ; n1059
g418 and n1050_not n1059 ; n1060
g419 and in2[76]_not in3[76] ; n1061
g420 and n722_not n1061_not ; n1062
g421 and n721 n1062 ; n1063
g422 and n1060_not n1063 ; n1064
g423 and n729_not n1064_not ; n1065
g424 and n727_not n1065 ; n1066
g425 and n718_not n1066 ; n1067
g426 and n717_not n1067_not ; n1068
g427 and n716 n1068 ; n1069
g428 and n713_not n1069 ; n1070
g429 and in2[83] in3[83]_not ; n1071
g430 and in3[80]_not n717_not ; n1072
g431 and in2[80] n1072 ; n1073
g432 and in2[81] in3[81]_not ; n1074
g433 and n1073_not n1074_not ; n1075
g434 and in2[82] in3[82]_not ; n1076
g435 and n1075 n1076_not ; n1077
g436 and n716 n1077_not ; n1078
g437 and n1071_not n1078_not ; n1079
g438 and n1070_not n1079 ; n1080
g439 and in2[84]_not in3[84] ; n1081
g440 and n705_not n1081_not ; n1082
g441 and n704 n1082 ; n1083
g442 and n1080_not n1083 ; n1084
g443 and n712_not n1084_not ; n1085
g444 and n710_not n1085 ; n1086
g445 and n701_not n1086 ; n1087
g446 and in2[91]_not in3[91] ; n1088
g447 and in2[90]_not in3[90] ; n1089
g448 and n1088_not n1089_not ; n1090
g449 and in2[89]_not in3[89] ; n1091
g450 and in2[88]_not in3[88] ; n1092
g451 and n1091_not n1092_not ; n1093
g452 and n1090 n1093 ; n1094
g453 and n1087_not n1094 ; n1095
g454 and in2[91] in3[91]_not ; n1096
g455 and in2[88] in3[88]_not ; n1097
g456 and n1091_not n1097 ; n1098
g457 and in2[89] in3[89]_not ; n1099
g458 and n1098_not n1099_not ; n1100
g459 and in2[90] in3[90]_not ; n1101
g460 and n1100 n1101_not ; n1102
g461 and n1090 n1102_not ; n1103
g462 and n1096_not n1103_not ; n1104
g463 and n1095_not n1104 ; n1105
g464 and in2[92]_not in3[92] ; n1106
g465 and n693_not n1106_not ; n1107
g466 and n692 n1107 ; n1108
g467 and n1105_not n1108 ; n1109
g468 and n700_not n1109_not ; n1110
g469 and n698_not n1110 ; n1111
g470 and n689_not n1111 ; n1112
g471 and n688_not n1112_not ; n1113
g472 and n687 n1113 ; n1114
g473 and n684_not n1114 ; n1115
g474 and in2[99] in3[99]_not ; n1116
g475 and in3[96]_not n688_not ; n1117
g476 and in2[96] n1117 ; n1118
g477 and in2[97] in3[97]_not ; n1119
g478 and n1118_not n1119_not ; n1120
g479 and in2[98] in3[98]_not ; n1121
g480 and n1120 n1121_not ; n1122
g481 and n687 n1122_not ; n1123
g482 and n1116_not n1123_not ; n1124
g483 and n1115_not n1124 ; n1125
g484 and in2[100]_not in3[100] ; n1126
g485 and n676_not n1126_not ; n1127
g486 and n675 n1127 ; n1128
g487 and n1125_not n1128 ; n1129
g488 and n683_not n1129_not ; n1130
g489 and n681_not n1130 ; n1131
g490 and n672_not n1131 ; n1132
g491 and in2[107]_not in3[107] ; n1133
g492 and in2[106]_not in3[106] ; n1134
g493 and n1133_not n1134_not ; n1135
g494 and in2[105]_not in3[105] ; n1136
g495 and in2[104]_not in3[104] ; n1137
g496 and n1136_not n1137_not ; n1138
g497 and n1135 n1138 ; n1139
g498 and n1132_not n1139 ; n1140
g499 and in2[107] in3[107]_not ; n1141
g500 and in2[104] in3[104]_not ; n1142
g501 and n1136_not n1142 ; n1143
g502 and in2[105] in3[105]_not ; n1144
g503 and n1143_not n1144_not ; n1145
g504 and in2[106] in3[106]_not ; n1146
g505 and n1145 n1146_not ; n1147
g506 and n1135 n1147_not ; n1148
g507 and n1141_not n1148_not ; n1149
g508 and n1140_not n1149 ; n1150
g509 and in2[108]_not in3[108] ; n1151
g510 and n664_not n1151_not ; n1152
g511 and n663 n1152 ; n1153
g512 and n1150_not n1153 ; n1154
g513 and n671_not n1154_not ; n1155
g514 and n669_not n1155 ; n1156
g515 and n660_not n1156 ; n1157
g516 and n659_not n1157_not ; n1158
g517 and n658 n1158 ; n1159
g518 and n655_not n1159 ; n1160
g519 and in2[115] in3[115]_not ; n1161
g520 and in3[112]_not n659_not ; n1162
g521 and in2[112] n1162 ; n1163
g522 and in2[113] in3[113]_not ; n1164
g523 and n1163_not n1164_not ; n1165
g524 and in2[114] in3[114]_not ; n1166
g525 and n1165 n1166_not ; n1167
g526 and n658 n1167_not ; n1168
g527 and n1161_not n1168_not ; n1169
g528 and n1160_not n1169 ; n1170
g529 and in2[116]_not in3[116] ; n1171
g530 and n647_not n1171_not ; n1172
g531 and n646 n1172 ; n1173
g532 and n1170_not n1173 ; n1174
g533 and n654_not n1174_not ; n1175
g534 and n652_not n1175 ; n1176
g535 and n643_not n1176 ; n1177
g536 and in2[123]_not in3[123] ; n1178
g537 and in2[122]_not in3[122] ; n1179
g538 and n1178_not n1179_not ; n1180
g539 and in2[121]_not in3[121] ; n1181
g540 and in2[120]_not in3[120] ; n1182
g541 and n1181_not n1182_not ; n1183
g542 and n1180 n1183 ; n1184
g543 and n1177_not n1184 ; n1185
g544 and in2[123] in3[123]_not ; n1186
g545 and in2[120] in3[120]_not ; n1187
g546 and n1181_not n1187 ; n1188
g547 and in2[121] in3[121]_not ; n1189
g548 and n1188_not n1189_not ; n1190
g549 and in2[122] in3[122]_not ; n1191
g550 and n1190 n1191_not ; n1192
g551 and n1180 n1192_not ; n1193
g552 and n1186_not n1193_not ; n1194
g553 and n1185_not n1194 ; n1195
g554 and in2[124]_not in3[124] ; n1196
g555 and in2[127] in3[127]_not ; n1197
g556 and in2[126]_not in3[126] ; n1198
g557 and in2[125]_not in3[125] ; n1199
g558 and n1198_not n1199_not ; n1200
g559 and n1197_not n1200 ; n1201
g560 and n1196_not n1201 ; n1202
g561 and n1195_not n1202 ; n1203
g562 and in2[124] in3[124]_not ; n1204
g563 and in2[125] in3[125]_not ; n1205
g564 and n1204_not n1205_not ; n1206
g565 and n1200 n1206_not ; n1207
g566 and in2[126] in3[126]_not ; n1208
g567 and n1207_not n1208_not ; n1209
g568 and n1197_not n1209_not ; n1210
g569 and n1203_not n1210_not ; n1211
g570 and in3[127]_not n1211 ; n1212
g571 and in2[127] n1212_not ; n1213
g572 and in0[119] in1[119]_not ; n1214
g573 and in0[119]_not in1[119] ; n1215
g574 and in0[118]_not in1[118] ; n1216
g575 and n1215_not n1216_not ; n1217
g576 and in0[117]_not in1[117] ; n1218
g577 and in0[116] in1[116]_not ; n1219
g578 and n1218_not n1219 ; n1220
g579 and in0[117] in1[117]_not ; n1221
g580 and n1220_not n1221_not ; n1222
g581 and n1217 n1222_not ; n1223
g582 and in1[118]_not n1215_not ; n1224
g583 and in0[118] n1224 ; n1225
g584 and in0[112]_not in1[112] ; n1226
g585 and in0[115]_not in1[115] ; n1227
g586 and in0[114]_not in1[114] ; n1228
g587 and n1227_not n1228_not ; n1229
g588 and in0[113]_not in1[113] ; n1230
g589 and in0[111] in1[111]_not ; n1231
g590 and in0[111]_not in1[111] ; n1232
g591 and in0[110]_not in1[110] ; n1233
g592 and n1232_not n1233_not ; n1234
g593 and in0[109]_not in1[109] ; n1235
g594 and in0[108] in1[108]_not ; n1236
g595 and n1235_not n1236 ; n1237
g596 and in0[109] in1[109]_not ; n1238
g597 and n1237_not n1238_not ; n1239
g598 and n1234 n1239_not ; n1240
g599 and in1[110]_not n1232_not ; n1241
g600 and in0[110] n1241 ; n1242
g601 and in0[103] in1[103]_not ; n1243
g602 and in0[103]_not in1[103] ; n1244
g603 and in0[102]_not in1[102] ; n1245
g604 and n1244_not n1245_not ; n1246
g605 and in0[101]_not in1[101] ; n1247
g606 and in0[100] in1[100]_not ; n1248
g607 and n1247_not n1248 ; n1249
g608 and in0[101] in1[101]_not ; n1250
g609 and n1249_not n1250_not ; n1251
g610 and n1246 n1251_not ; n1252
g611 and in1[102]_not n1244_not ; n1253
g612 and in0[102] n1253 ; n1254
g613 and in0[96]_not in1[96] ; n1255
g614 and in0[99]_not in1[99] ; n1256
g615 and in0[98]_not in1[98] ; n1257
g616 and n1256_not n1257_not ; n1258
g617 and in0[97]_not in1[97] ; n1259
g618 and in0[95] in1[95]_not ; n1260
g619 and in0[95]_not in1[95] ; n1261
g620 and in0[94]_not in1[94] ; n1262
g621 and n1261_not n1262_not ; n1263
g622 and in0[93]_not in1[93] ; n1264
g623 and in0[92] in1[92]_not ; n1265
g624 and n1264_not n1265 ; n1266
g625 and in0[93] in1[93]_not ; n1267
g626 and n1266_not n1267_not ; n1268
g627 and n1263 n1268_not ; n1269
g628 and in1[94]_not n1261_not ; n1270
g629 and in0[94] n1270 ; n1271
g630 and in0[87] in1[87]_not ; n1272
g631 and in0[87]_not in1[87] ; n1273
g632 and in0[86]_not in1[86] ; n1274
g633 and n1273_not n1274_not ; n1275
g634 and in0[85]_not in1[85] ; n1276
g635 and in0[84] in1[84]_not ; n1277
g636 and n1276_not n1277 ; n1278
g637 and in0[85] in1[85]_not ; n1279
g638 and n1278_not n1279_not ; n1280
g639 and n1275 n1280_not ; n1281
g640 and in1[86]_not n1273_not ; n1282
g641 and in0[86] n1282 ; n1283
g642 and in0[80]_not in1[80] ; n1284
g643 and in0[83]_not in1[83] ; n1285
g644 and in0[82]_not in1[82] ; n1286
g645 and n1285_not n1286_not ; n1287
g646 and in0[81]_not in1[81] ; n1288
g647 and in0[79] in1[79]_not ; n1289
g648 and in0[79]_not in1[79] ; n1290
g649 and in0[78]_not in1[78] ; n1291
g650 and n1290_not n1291_not ; n1292
g651 and in0[77]_not in1[77] ; n1293
g652 and in0[76] in1[76]_not ; n1294
g653 and n1293_not n1294 ; n1295
g654 and in0[77] in1[77]_not ; n1296
g655 and n1295_not n1296_not ; n1297
g656 and n1292 n1297_not ; n1298
g657 and in1[78]_not n1290_not ; n1299
g658 and in0[78] n1299 ; n1300
g659 and in0[71] in1[71]_not ; n1301
g660 and in0[71]_not in1[71] ; n1302
g661 and in0[70]_not in1[70] ; n1303
g662 and n1302_not n1303_not ; n1304
g663 and in0[69]_not in1[69] ; n1305
g664 and in0[68] in1[68]_not ; n1306
g665 and n1305_not n1306 ; n1307
g666 and in0[69] in1[69]_not ; n1308
g667 and n1307_not n1308_not ; n1309
g668 and n1304 n1309_not ; n1310
g669 and in1[70]_not n1302_not ; n1311
g670 and in0[70] n1311 ; n1312
g671 and in0[67]_not in1[67] ; n1313
g672 and in0[66]_not in1[66] ; n1314
g673 and n1313_not n1314_not ; n1315
g674 and in0[65]_not in1[65] ; n1316
g675 and in0[63] in1[63]_not ; n1317
g676 and in0[63]_not in1[63] ; n1318
g677 and in0[62]_not in1[62] ; n1319
g678 and n1318_not n1319_not ; n1320
g679 and in0[60]_not in1[60] ; n1321
g680 and in0[61]_not in1[61] ; n1322
g681 and n1321_not n1322_not ; n1323
g682 and n1320 n1323 ; n1324
g683 and in0[59] in1[59]_not ; n1325
g684 and in0[59]_not in1[59] ; n1326
g685 and in0[58]_not in1[58] ; n1327
g686 and n1326_not n1327_not ; n1328
g687 and in0[57]_not in1[57] ; n1329
g688 and in0[56] in1[56]_not ; n1330
g689 and n1329_not n1330 ; n1331
g690 and in0[57] in1[57]_not ; n1332
g691 and n1331_not n1332_not ; n1333
g692 and in0[58] in1[58]_not ; n1334
g693 and n1333 n1334_not ; n1335
g694 and n1328 n1335_not ; n1336
g695 and n1325_not n1336_not ; n1337
g696 and n1324 n1337_not ; n1338
g697 and in0[60] in1[60]_not ; n1339
g698 and n1322_not n1339 ; n1340
g699 and in0[61] in1[61]_not ; n1341
g700 and n1340_not n1341_not ; n1342
g701 and n1320 n1342_not ; n1343
g702 and in1[62]_not n1318_not ; n1344
g703 and in0[62] n1344 ; n1345
g704 and in0[47] in1[47]_not ; n1346
g705 and in0[47]_not in1[47] ; n1347
g706 and in0[46]_not in1[46] ; n1348
g707 and n1347_not n1348_not ; n1349
g708 and in0[44]_not in1[44] ; n1350
g709 and in0[45]_not in1[45] ; n1351
g710 and n1350_not n1351_not ; n1352
g711 and n1349 n1352 ; n1353
g712 and in0[43] in1[43]_not ; n1354
g713 and in0[43]_not in1[43] ; n1355
g714 and in0[42]_not in1[42] ; n1356
g715 and n1355_not n1356_not ; n1357
g716 and in0[41]_not in1[41] ; n1358
g717 and in0[40] in1[40]_not ; n1359
g718 and n1358_not n1359 ; n1360
g719 and in0[41] in1[41]_not ; n1361
g720 and n1360_not n1361_not ; n1362
g721 and in0[42] in1[42]_not ; n1363
g722 and n1362 n1363_not ; n1364
g723 and n1357 n1364_not ; n1365
g724 and n1354_not n1365_not ; n1366
g725 and n1353 n1366_not ; n1367
g726 and in0[44] in1[44]_not ; n1368
g727 and n1351_not n1368 ; n1369
g728 and in0[45] in1[45]_not ; n1370
g729 and n1369_not n1370_not ; n1371
g730 and n1349 n1371_not ; n1372
g731 and in1[46]_not n1347_not ; n1373
g732 and in0[46] n1373 ; n1374
g733 and in0[32]_not in1[32] ; n1375
g734 and in0[31]_not in1[31] ; n1376
g735 and in0[30]_not in1[30] ; n1377
g736 and in0[29]_not in1[29] ; n1378
g737 and in0[28]_not in1[28] ; n1379
g738 and in0[27]_not in1[27] ; n1380
g739 and in0[26]_not in1[26] ; n1381
g740 and in0[23]_not in1[23] ; n1382
g741 and in0[22]_not in1[22] ; n1383
g742 and in0[21]_not in1[21] ; n1384
g743 and in0[20]_not in1[20] ; n1385
g744 and in0[19]_not in1[19] ; n1386
g745 and in0[18]_not in1[18] ; n1387
g746 and in0[15]_not in1[15] ; n1388
g747 and in0[14]_not in1[14] ; n1389
g748 and in0[13]_not in1[13] ; n1390
g749 and in0[12]_not in1[12] ; n1391
g750 and in0[11]_not in1[11] ; n1392
g751 and in0[10]_not in1[10] ; n1393
g752 and in0[7]_not in1[7] ; n1394
g753 and in0[6]_not in1[6] ; n1395
g754 and in0[3]_not in1[3] ; n1396
g755 and in0[0] in1[0]_not ; n1397
g756 and in0[1] in1[1]_not ; n1398
g757 and n1397_not n1398_not ; n1399
g758 and in0[2]_not in1[2] ; n1400
g759 and in0[1]_not in1[1] ; n1401
g760 and n1400_not n1401_not ; n1402
g761 and n1399_not n1402 ; n1403
g762 and in0[2] in1[2]_not ; n1404
g763 and n1403_not n1404_not ; n1405
g764 and n1396_not n1405_not ; n1406
g765 and in0[3] in1[3]_not ; n1407
g766 and n1406_not n1407_not ; n1408
g767 and in0[4]_not n1408 ; n1409
g768 and in1[4]_not n1409_not ; n1410
g769 and in0[4] n1408_not ; n1411
g770 and n1410_not n1411_not ; n1412
g771 and in0[5]_not n1412 ; n1413
g772 and in1[5]_not n1413_not ; n1414
g773 and in0[5] n1412_not ; n1415
g774 and n1414_not n1415_not ; n1416
g775 and n1395_not n1416_not ; n1417
g776 and in0[6] in1[6]_not ; n1418
g777 and n1417_not n1418_not ; n1419
g778 and n1394_not n1419_not ; n1420
g779 and in0[7] in1[7]_not ; n1421
g780 and n1420_not n1421_not ; n1422
g781 and in0[8]_not n1422 ; n1423
g782 and in1[8]_not n1423_not ; n1424
g783 and in0[8] n1422_not ; n1425
g784 and n1424_not n1425_not ; n1426
g785 and in0[9]_not n1426 ; n1427
g786 and in1[9]_not n1427_not ; n1428
g787 and in0[9] n1426_not ; n1429
g788 and n1428_not n1429_not ; n1430
g789 and n1393_not n1430_not ; n1431
g790 and in0[10] in1[10]_not ; n1432
g791 and n1431_not n1432_not ; n1433
g792 and n1392_not n1433_not ; n1434
g793 and in0[11] in1[11]_not ; n1435
g794 and n1434_not n1435_not ; n1436
g795 and n1391_not n1436_not ; n1437
g796 and in0[12] in1[12]_not ; n1438
g797 and n1437_not n1438_not ; n1439
g798 and n1390_not n1439_not ; n1440
g799 and in0[13] in1[13]_not ; n1441
g800 and n1440_not n1441_not ; n1442
g801 and n1389_not n1442_not ; n1443
g802 and in0[14] in1[14]_not ; n1444
g803 and n1443_not n1444_not ; n1445
g804 and n1388_not n1445_not ; n1446
g805 and in0[15] in1[15]_not ; n1447
g806 and n1446_not n1447_not ; n1448
g807 and in0[16]_not n1448 ; n1449
g808 and in1[16]_not n1449_not ; n1450
g809 and in0[16] n1448_not ; n1451
g810 and n1450_not n1451_not ; n1452
g811 and in0[17]_not n1452 ; n1453
g812 and in1[17]_not n1453_not ; n1454
g813 and in0[17] n1452_not ; n1455
g814 and n1454_not n1455_not ; n1456
g815 and n1387_not n1456_not ; n1457
g816 and in0[18] in1[18]_not ; n1458
g817 and n1457_not n1458_not ; n1459
g818 and n1386_not n1459_not ; n1460
g819 and in0[19] in1[19]_not ; n1461
g820 and n1460_not n1461_not ; n1462
g821 and n1385_not n1462_not ; n1463
g822 and in0[20] in1[20]_not ; n1464
g823 and n1463_not n1464_not ; n1465
g824 and n1384_not n1465_not ; n1466
g825 and in0[21] in1[21]_not ; n1467
g826 and n1466_not n1467_not ; n1468
g827 and n1383_not n1468_not ; n1469
g828 and in0[22] in1[22]_not ; n1470
g829 and n1469_not n1470_not ; n1471
g830 and n1382_not n1471_not ; n1472
g831 and in0[23] in1[23]_not ; n1473
g832 and n1472_not n1473_not ; n1474
g833 and in0[24]_not n1474 ; n1475
g834 and in1[24]_not n1475_not ; n1476
g835 and in0[24] n1474_not ; n1477
g836 and n1476_not n1477_not ; n1478
g837 and in0[25]_not n1478 ; n1479
g838 and in1[25]_not n1479_not ; n1480
g839 and in0[25] n1478_not ; n1481
g840 and n1480_not n1481_not ; n1482
g841 and n1381_not n1482_not ; n1483
g842 and in0[26] in1[26]_not ; n1484
g843 and n1483_not n1484_not ; n1485
g844 and n1380_not n1485_not ; n1486
g845 and in0[27] in1[27]_not ; n1487
g846 and n1486_not n1487_not ; n1488
g847 and n1379_not n1488_not ; n1489
g848 and in0[28] in1[28]_not ; n1490
g849 and n1489_not n1490_not ; n1491
g850 and n1378_not n1491_not ; n1492
g851 and in0[29] in1[29]_not ; n1493
g852 and n1492_not n1493_not ; n1494
g853 and n1377_not n1494_not ; n1495
g854 and in0[30] in1[30]_not ; n1496
g855 and n1495_not n1496_not ; n1497
g856 and n1376_not n1497_not ; n1498
g857 and in0[31] in1[31]_not ; n1499
g858 and n1498_not n1499_not ; n1500
g859 and in0[39]_not in1[39] ; n1501
g860 and in0[38]_not in1[38] ; n1502
g861 and n1501_not n1502_not ; n1503
g862 and in0[36]_not in1[36] ; n1504
g863 and in0[37]_not in1[37] ; n1505
g864 and n1504_not n1505_not ; n1506
g865 and n1503 n1506 ; n1507
g866 and in0[33]_not in1[33] ; n1508
g867 and in0[35]_not in1[35] ; n1509
g868 and in0[34]_not in1[34] ; n1510
g869 and n1509_not n1510_not ; n1511
g870 and n1508_not n1511 ; n1512
g871 and n1507 n1512 ; n1513
g872 and n1500_not n1513 ; n1514
g873 and n1375_not n1514 ; n1515
g874 and in0[39] in1[39]_not ; n1516
g875 and in0[36] in1[36]_not ; n1517
g876 and n1505_not n1517 ; n1518
g877 and in0[37] in1[37]_not ; n1519
g878 and n1518_not n1519_not ; n1520
g879 and n1503 n1520_not ; n1521
g880 and in1[38]_not n1501_not ; n1522
g881 and in0[38] n1522 ; n1523
g882 and in0[35] in1[35]_not ; n1524
g883 and in1[32]_not n1508_not ; n1525
g884 and in0[32] n1525 ; n1526
g885 and in0[33] in1[33]_not ; n1527
g886 and n1526_not n1527_not ; n1528
g887 and in0[34] in1[34]_not ; n1529
g888 and n1528 n1529_not ; n1530
g889 and n1511 n1530_not ; n1531
g890 and n1524_not n1531_not ; n1532
g891 and n1507 n1532_not ; n1533
g892 and n1523_not n1533_not ; n1534
g893 and n1521_not n1534 ; n1535
g894 and n1516_not n1535 ; n1536
g895 and n1515_not n1536 ; n1537
g896 and in0[40]_not in1[40] ; n1538
g897 and n1358_not n1538_not ; n1539
g898 and n1357 n1539 ; n1540
g899 and n1353 n1540 ; n1541
g900 and n1537_not n1541 ; n1542
g901 and n1374_not n1542_not ; n1543
g902 and n1372_not n1543 ; n1544
g903 and n1367_not n1544 ; n1545
g904 and n1346_not n1545 ; n1546
g905 and in0[48]_not in1[48] ; n1547
g906 and in0[55]_not in1[55] ; n1548
g907 and in0[54]_not in1[54] ; n1549
g908 and n1548_not n1549_not ; n1550
g909 and in0[53]_not in1[53] ; n1551
g910 and in0[52]_not in1[52] ; n1552
g911 and n1551_not n1552_not ; n1553
g912 and n1550 n1553 ; n1554
g913 and in0[49]_not in1[49] ; n1555
g914 and in0[51]_not in1[51] ; n1556
g915 and in0[50]_not in1[50] ; n1557
g916 and n1556_not n1557_not ; n1558
g917 and n1555_not n1558 ; n1559
g918 and n1554 n1559 ; n1560
g919 and n1547_not n1560 ; n1561
g920 and n1546_not n1561 ; n1562
g921 and in0[55] in1[55]_not ; n1563
g922 and in0[51] in1[51]_not ; n1564
g923 and in1[48]_not n1555_not ; n1565
g924 and in0[48] n1565 ; n1566
g925 and in0[49] in1[49]_not ; n1567
g926 and n1566_not n1567_not ; n1568
g927 and in0[50] in1[50]_not ; n1569
g928 and n1568 n1569_not ; n1570
g929 and n1558 n1570_not ; n1571
g930 and n1564_not n1571_not ; n1572
g931 and n1554 n1572_not ; n1573
g932 and in0[52] in1[52]_not ; n1574
g933 and n1551_not n1574 ; n1575
g934 and in0[53] in1[53]_not ; n1576
g935 and n1575_not n1576_not ; n1577
g936 and in0[54] in1[54]_not ; n1578
g937 and n1577 n1578_not ; n1579
g938 and n1550 n1579_not ; n1580
g939 and n1573_not n1580_not ; n1581
g940 and n1563_not n1581 ; n1582
g941 and n1562_not n1582 ; n1583
g942 and in0[56]_not in1[56] ; n1584
g943 and n1329_not n1584_not ; n1585
g944 and n1324 n1585 ; n1586
g945 and n1328 n1586 ; n1587
g946 and n1583_not n1587 ; n1588
g947 and n1345_not n1588_not ; n1589
g948 and n1343_not n1589 ; n1590
g949 and n1338_not n1590 ; n1591
g950 and n1317_not n1591 ; n1592
g951 and in0[64]_not in1[64] ; n1593
g952 and n1592_not n1593_not ; n1594
g953 and n1316_not n1594 ; n1595
g954 and n1315 n1595 ; n1596
g955 and in0[67] in1[67]_not ; n1597
g956 and in0[64] in1[64]_not ; n1598
g957 and n1316_not n1598 ; n1599
g958 and in0[65] in1[65]_not ; n1600
g959 and n1599_not n1600_not ; n1601
g960 and in0[66] in1[66]_not ; n1602
g961 and n1601 n1602_not ; n1603
g962 and n1315 n1603_not ; n1604
g963 and n1597_not n1604_not ; n1605
g964 and n1596_not n1605 ; n1606
g965 and in0[68]_not in1[68] ; n1607
g966 and n1305_not n1607_not ; n1608
g967 and n1304 n1608 ; n1609
g968 and n1606_not n1609 ; n1610
g969 and n1312_not n1610_not ; n1611
g970 and n1310_not n1611 ; n1612
g971 and n1301_not n1612 ; n1613
g972 and in0[75]_not in1[75] ; n1614
g973 and in0[74]_not in1[74] ; n1615
g974 and n1614_not n1615_not ; n1616
g975 and in0[73]_not in1[73] ; n1617
g976 and in0[72]_not in1[72] ; n1618
g977 and n1617_not n1618_not ; n1619
g978 and n1616 n1619 ; n1620
g979 and n1613_not n1620 ; n1621
g980 and in0[75] in1[75]_not ; n1622
g981 and in0[72] in1[72]_not ; n1623
g982 and n1617_not n1623 ; n1624
g983 and in0[73] in1[73]_not ; n1625
g984 and n1624_not n1625_not ; n1626
g985 and in0[74] in1[74]_not ; n1627
g986 and n1626 n1627_not ; n1628
g987 and n1616 n1628_not ; n1629
g988 and n1622_not n1629_not ; n1630
g989 and n1621_not n1630 ; n1631
g990 and in0[76]_not in1[76] ; n1632
g991 and n1293_not n1632_not ; n1633
g992 and n1292 n1633 ; n1634
g993 and n1631_not n1634 ; n1635
g994 and n1300_not n1635_not ; n1636
g995 and n1298_not n1636 ; n1637
g996 and n1289_not n1637 ; n1638
g997 and n1288_not n1638_not ; n1639
g998 and n1287 n1639 ; n1640
g999 and n1284_not n1640 ; n1641
g1000 and in0[83] in1[83]_not ; n1642
g1001 and in1[80]_not n1288_not ; n1643
g1002 and in0[80] n1643 ; n1644
g1003 and in0[81] in1[81]_not ; n1645
g1004 and n1644_not n1645_not ; n1646
g1005 and in0[82] in1[82]_not ; n1647
g1006 and n1646 n1647_not ; n1648
g1007 and n1287 n1648_not ; n1649
g1008 and n1642_not n1649_not ; n1650
g1009 and n1641_not n1650 ; n1651
g1010 and in0[84]_not in1[84] ; n1652
g1011 and n1276_not n1652_not ; n1653
g1012 and n1275 n1653 ; n1654
g1013 and n1651_not n1654 ; n1655
g1014 and n1283_not n1655_not ; n1656
g1015 and n1281_not n1656 ; n1657
g1016 and n1272_not n1657 ; n1658
g1017 and in0[91]_not in1[91] ; n1659
g1018 and in0[90]_not in1[90] ; n1660
g1019 and n1659_not n1660_not ; n1661
g1020 and in0[89]_not in1[89] ; n1662
g1021 and in0[88]_not in1[88] ; n1663
g1022 and n1662_not n1663_not ; n1664
g1023 and n1661 n1664 ; n1665
g1024 and n1658_not n1665 ; n1666
g1025 and in0[91] in1[91]_not ; n1667
g1026 and in0[88] in1[88]_not ; n1668
g1027 and n1662_not n1668 ; n1669
g1028 and in0[89] in1[89]_not ; n1670
g1029 and n1669_not n1670_not ; n1671
g1030 and in0[90] in1[90]_not ; n1672
g1031 and n1671 n1672_not ; n1673
g1032 and n1661 n1673_not ; n1674
g1033 and n1667_not n1674_not ; n1675
g1034 and n1666_not n1675 ; n1676
g1035 and in0[92]_not in1[92] ; n1677
g1036 and n1264_not n1677_not ; n1678
g1037 and n1263 n1678 ; n1679
g1038 and n1676_not n1679 ; n1680
g1039 and n1271_not n1680_not ; n1681
g1040 and n1269_not n1681 ; n1682
g1041 and n1260_not n1682 ; n1683
g1042 and n1259_not n1683_not ; n1684
g1043 and n1258 n1684 ; n1685
g1044 and n1255_not n1685 ; n1686
g1045 and in0[99] in1[99]_not ; n1687
g1046 and in1[96]_not n1259_not ; n1688
g1047 and in0[96] n1688 ; n1689
g1048 and in0[97] in1[97]_not ; n1690
g1049 and n1689_not n1690_not ; n1691
g1050 and in0[98] in1[98]_not ; n1692
g1051 and n1691 n1692_not ; n1693
g1052 and n1258 n1693_not ; n1694
g1053 and n1687_not n1694_not ; n1695
g1054 and n1686_not n1695 ; n1696
g1055 and in0[100]_not in1[100] ; n1697
g1056 and n1247_not n1697_not ; n1698
g1057 and n1246 n1698 ; n1699
g1058 and n1696_not n1699 ; n1700
g1059 and n1254_not n1700_not ; n1701
g1060 and n1252_not n1701 ; n1702
g1061 and n1243_not n1702 ; n1703
g1062 and in0[107]_not in1[107] ; n1704
g1063 and in0[106]_not in1[106] ; n1705
g1064 and n1704_not n1705_not ; n1706
g1065 and in0[105]_not in1[105] ; n1707
g1066 and in0[104]_not in1[104] ; n1708
g1067 and n1707_not n1708_not ; n1709
g1068 and n1706 n1709 ; n1710
g1069 and n1703_not n1710 ; n1711
g1070 and in0[107] in1[107]_not ; n1712
g1071 and in0[104] in1[104]_not ; n1713
g1072 and n1707_not n1713 ; n1714
g1073 and in0[105] in1[105]_not ; n1715
g1074 and n1714_not n1715_not ; n1716
g1075 and in0[106] in1[106]_not ; n1717
g1076 and n1716 n1717_not ; n1718
g1077 and n1706 n1718_not ; n1719
g1078 and n1712_not n1719_not ; n1720
g1079 and n1711_not n1720 ; n1721
g1080 and in0[108]_not in1[108] ; n1722
g1081 and n1235_not n1722_not ; n1723
g1082 and n1234 n1723 ; n1724
g1083 and n1721_not n1724 ; n1725
g1084 and n1242_not n1725_not ; n1726
g1085 and n1240_not n1726 ; n1727
g1086 and n1231_not n1727 ; n1728
g1087 and n1230_not n1728_not ; n1729
g1088 and n1229 n1729 ; n1730
g1089 and n1226_not n1730 ; n1731
g1090 and in0[115] in1[115]_not ; n1732
g1091 and in1[112]_not n1230_not ; n1733
g1092 and in0[112] n1733 ; n1734
g1093 and in0[113] in1[113]_not ; n1735
g1094 and n1734_not n1735_not ; n1736
g1095 and in0[114] in1[114]_not ; n1737
g1096 and n1736 n1737_not ; n1738
g1097 and n1229 n1738_not ; n1739
g1098 and n1732_not n1739_not ; n1740
g1099 and n1731_not n1740 ; n1741
g1100 and in0[116]_not in1[116] ; n1742
g1101 and n1218_not n1742_not ; n1743
g1102 and n1217 n1743 ; n1744
g1103 and n1741_not n1744 ; n1745
g1104 and n1225_not n1745_not ; n1746
g1105 and n1223_not n1746 ; n1747
g1106 and n1214_not n1747 ; n1748
g1107 and in0[123]_not in1[123] ; n1749
g1108 and in0[122]_not in1[122] ; n1750
g1109 and n1749_not n1750_not ; n1751
g1110 and in0[121]_not in1[121] ; n1752
g1111 and in0[120]_not in1[120] ; n1753
g1112 and n1752_not n1753_not ; n1754
g1113 and n1751 n1754 ; n1755
g1114 and n1748_not n1755 ; n1756
g1115 and in0[123] in1[123]_not ; n1757
g1116 and in0[120] in1[120]_not ; n1758
g1117 and n1752_not n1758 ; n1759
g1118 and in0[121] in1[121]_not ; n1760
g1119 and n1759_not n1760_not ; n1761
g1120 and in0[122] in1[122]_not ; n1762
g1121 and n1761 n1762_not ; n1763
g1122 and n1751 n1763_not ; n1764
g1123 and n1757_not n1764_not ; n1765
g1124 and n1756_not n1765 ; n1766
g1125 and in0[124]_not in1[124] ; n1767
g1126 and in0[127] in1[127]_not ; n1768
g1127 and in0[126]_not in1[126] ; n1769
g1128 and in0[125]_not in1[125] ; n1770
g1129 and n1769_not n1770_not ; n1771
g1130 and n1768_not n1771 ; n1772
g1131 and n1767_not n1772 ; n1773
g1132 and n1766_not n1773 ; n1774
g1133 and in0[124] in1[124]_not ; n1775
g1134 and in0[125] in1[125]_not ; n1776
g1135 and n1775_not n1776_not ; n1777
g1136 and n1771 n1777_not ; n1778
g1137 and in0[126] in1[126]_not ; n1779
g1138 and n1778_not n1779_not ; n1780
g1139 and n1768_not n1780_not ; n1781
g1140 and n1774_not n1781_not ; n1782
g1141 and in1[127]_not n1782 ; n1783
g1142 and in0[127] n1783_not ; n1784
g1143 and n1213 n1784_not ; n1785
g1144 and in0[127]_not in1[127] ; n1786
g1145 and n1782 n1786_not ; n1787
g1146 and in1[119] n1787 ; n1788
g1147 and in0[119] n1787_not ; n1789
g1148 and n1788_not n1789_not ; n1790
g1149 and in2[127]_not in3[127] ; n1791
g1150 and n1211 n1791_not ; n1792
g1151 and in3[119] n1792 ; n1793
g1152 and in2[119] n1792_not ; n1794
g1153 and n1793_not n1794_not ; n1795
g1154 and n1790_not n1795 ; n1796
g1155 and n1790 n1795_not ; n1797
g1156 and in3[118] n1792 ; n1798
g1157 and in2[118] n1792_not ; n1799
g1158 and n1798_not n1799_not ; n1800
g1159 and in1[118] n1787 ; n1801
g1160 and in0[118] n1787_not ; n1802
g1161 and n1801_not n1802_not ; n1803
g1162 and n1800_not n1803 ; n1804
g1163 and n1797_not n1804_not ; n1805
g1164 and in1[116] n1787 ; n1806
g1165 and in0[116] n1787_not ; n1807
g1166 and n1806_not n1807_not ; n1808
g1167 and in1[117] n1787 ; n1809
g1168 and in0[117] n1787_not ; n1810
g1169 and n1809_not n1810_not ; n1811
g1170 and in3[117] n1792 ; n1812
g1171 and in2[117] n1792_not ; n1813
g1172 and n1812_not n1813_not ; n1814
g1173 and n1811 n1814_not ; n1815
g1174 and in3[116] n1792 ; n1816
g1175 and in2[116] n1792_not ; n1817
g1176 and n1816_not n1817_not ; n1818
g1177 and n1815_not n1818 ; n1819
g1178 and n1808_not n1819 ; n1820
g1179 and n1811_not n1814 ; n1821
g1180 and n1820_not n1821_not ; n1822
g1181 and n1805 n1822_not ; n1823
g1182 and n1800 n1803_not ; n1824
g1183 and n1797_not n1824 ; n1825
g1184 and in3[112] n1792 ; n1826
g1185 and in2[112] n1792_not ; n1827
g1186 and n1826_not n1827_not ; n1828
g1187 and in1[112] n1787 ; n1829
g1188 and in0[112] n1787_not ; n1830
g1189 and n1829_not n1830_not ; n1831
g1190 and n1828_not n1831 ; n1832
g1191 and in1[115] n1787 ; n1833
g1192 and in0[115] n1787_not ; n1834
g1193 and n1833_not n1834_not ; n1835
g1194 and in3[115] n1792 ; n1836
g1195 and in2[115] n1792_not ; n1837
g1196 and n1836_not n1837_not ; n1838
g1197 and n1835 n1838_not ; n1839
g1198 and in3[114] n1792 ; n1840
g1199 and in2[114] n1792_not ; n1841
g1200 and n1840_not n1841_not ; n1842
g1201 and in1[114] n1787 ; n1843
g1202 and in0[114] n1787_not ; n1844
g1203 and n1843_not n1844_not ; n1845
g1204 and n1842_not n1845 ; n1846
g1205 and n1839_not n1846_not ; n1847
g1206 and in1[113] n1787 ; n1848
g1207 and in0[113] n1787_not ; n1849
g1208 and n1848_not n1849_not ; n1850
g1209 and in3[113] n1792 ; n1851
g1210 and in2[113] n1792_not ; n1852
g1211 and n1851_not n1852_not ; n1853
g1212 and n1850 n1853_not ; n1854
g1213 and in1[111] n1787 ; n1855
g1214 and in0[111] n1787_not ; n1856
g1215 and n1855_not n1856_not ; n1857
g1216 and in3[111] n1792 ; n1858
g1217 and in2[111] n1792_not ; n1859
g1218 and n1858_not n1859_not ; n1860
g1219 and n1857_not n1860 ; n1861
g1220 and n1857 n1860_not ; n1862
g1221 and in3[110] n1792 ; n1863
g1222 and in2[110] n1792_not ; n1864
g1223 and n1863_not n1864_not ; n1865
g1224 and in1[110] n1787 ; n1866
g1225 and in0[110] n1787_not ; n1867
g1226 and n1866_not n1867_not ; n1868
g1227 and n1865_not n1868 ; n1869
g1228 and n1862_not n1869_not ; n1870
g1229 and in1[109] n1787 ; n1871
g1230 and in0[109] n1787_not ; n1872
g1231 and n1871_not n1872_not ; n1873
g1232 and in3[109] n1792 ; n1874
g1233 and in2[109] n1792_not ; n1875
g1234 and n1874_not n1875_not ; n1876
g1235 and n1873 n1876_not ; n1877
g1236 and in1[108] n1787 ; n1878
g1237 and in0[108] n1787_not ; n1879
g1238 and n1878_not n1879_not ; n1880
g1239 and in3[108] n1792 ; n1881
g1240 and in2[108] n1792_not ; n1882
g1241 and n1881_not n1882_not ; n1883
g1242 and n1880_not n1883 ; n1884
g1243 and n1877_not n1884 ; n1885
g1244 and n1873_not n1876 ; n1886
g1245 and n1885_not n1886_not ; n1887
g1246 and n1870 n1887_not ; n1888
g1247 and n1865 n1868_not ; n1889
g1248 and n1862_not n1889 ; n1890
g1249 and in1[103] n1787 ; n1891
g1250 and in0[103] n1787_not ; n1892
g1251 and n1891_not n1892_not ; n1893
g1252 and in3[103] n1792 ; n1894
g1253 and in2[103] n1792_not ; n1895
g1254 and n1894_not n1895_not ; n1896
g1255 and n1893_not n1896 ; n1897
g1256 and n1893 n1896_not ; n1898
g1257 and in3[102] n1792 ; n1899
g1258 and in2[102] n1792_not ; n1900
g1259 and n1899_not n1900_not ; n1901
g1260 and in1[102] n1787 ; n1902
g1261 and in0[102] n1787_not ; n1903
g1262 and n1902_not n1903_not ; n1904
g1263 and n1901_not n1904 ; n1905
g1264 and n1898_not n1905_not ; n1906
g1265 and in1[101] n1787 ; n1907
g1266 and in0[101] n1787_not ; n1908
g1267 and n1907_not n1908_not ; n1909
g1268 and in3[101] n1792 ; n1910
g1269 and in2[101] n1792_not ; n1911
g1270 and n1910_not n1911_not ; n1912
g1271 and n1909 n1912_not ; n1913
g1272 and in1[100] n1787 ; n1914
g1273 and in0[100] n1787_not ; n1915
g1274 and n1914_not n1915_not ; n1916
g1275 and in3[100] n1792 ; n1917
g1276 and in2[100] n1792_not ; n1918
g1277 and n1917_not n1918_not ; n1919
g1278 and n1916_not n1919 ; n1920
g1279 and n1913_not n1920 ; n1921
g1280 and n1909_not n1912 ; n1922
g1281 and n1921_not n1922_not ; n1923
g1282 and n1906 n1923_not ; n1924
g1283 and n1901 n1904_not ; n1925
g1284 and n1898_not n1925 ; n1926
g1285 and in3[96] n1792 ; n1927
g1286 and in2[96] n1792_not ; n1928
g1287 and n1927_not n1928_not ; n1929
g1288 and in1[96] n1787 ; n1930
g1289 and in0[96] n1787_not ; n1931
g1290 and n1930_not n1931_not ; n1932
g1291 and n1929_not n1932 ; n1933
g1292 and in1[99] n1787 ; n1934
g1293 and in0[99] n1787_not ; n1935
g1294 and n1934_not n1935_not ; n1936
g1295 and in3[99] n1792 ; n1937
g1296 and in2[99] n1792_not ; n1938
g1297 and n1937_not n1938_not ; n1939
g1298 and n1936 n1939_not ; n1940
g1299 and in3[98] n1792 ; n1941
g1300 and in2[98] n1792_not ; n1942
g1301 and n1941_not n1942_not ; n1943
g1302 and in1[98] n1787 ; n1944
g1303 and in0[98] n1787_not ; n1945
g1304 and n1944_not n1945_not ; n1946
g1305 and n1943_not n1946 ; n1947
g1306 and n1940_not n1947_not ; n1948
g1307 and in1[97] n1787 ; n1949
g1308 and in0[97] n1787_not ; n1950
g1309 and n1949_not n1950_not ; n1951
g1310 and in3[97] n1792 ; n1952
g1311 and in2[97] n1792_not ; n1953
g1312 and n1952_not n1953_not ; n1954
g1313 and n1951 n1954_not ; n1955
g1314 and in1[95] n1787 ; n1956
g1315 and in0[95] n1787_not ; n1957
g1316 and n1956_not n1957_not ; n1958
g1317 and in3[95] n1792 ; n1959
g1318 and in2[95] n1792_not ; n1960
g1319 and n1959_not n1960_not ; n1961
g1320 and n1958_not n1961 ; n1962
g1321 and n1958 n1961_not ; n1963
g1322 and in3[94] n1792 ; n1964
g1323 and in2[94] n1792_not ; n1965
g1324 and n1964_not n1965_not ; n1966
g1325 and in1[94] n1787 ; n1967
g1326 and in0[94] n1787_not ; n1968
g1327 and n1967_not n1968_not ; n1969
g1328 and n1966_not n1969 ; n1970
g1329 and n1963_not n1970_not ; n1971
g1330 and in1[93] n1787 ; n1972
g1331 and in0[93] n1787_not ; n1973
g1332 and n1972_not n1973_not ; n1974
g1333 and in3[93] n1792 ; n1975
g1334 and in2[93] n1792_not ; n1976
g1335 and n1975_not n1976_not ; n1977
g1336 and n1974 n1977_not ; n1978
g1337 and in1[92] n1787 ; n1979
g1338 and in0[92] n1787_not ; n1980
g1339 and n1979_not n1980_not ; n1981
g1340 and in3[92] n1792 ; n1982
g1341 and in2[92] n1792_not ; n1983
g1342 and n1982_not n1983_not ; n1984
g1343 and n1981_not n1984 ; n1985
g1344 and n1978_not n1985 ; n1986
g1345 and n1974_not n1977 ; n1987
g1346 and n1986_not n1987_not ; n1988
g1347 and n1971 n1988_not ; n1989
g1348 and n1966 n1969_not ; n1990
g1349 and n1963_not n1990 ; n1991
g1350 and in1[87] n1787 ; n1992
g1351 and in0[87] n1787_not ; n1993
g1352 and n1992_not n1993_not ; n1994
g1353 and in3[87] n1792 ; n1995
g1354 and in2[87] n1792_not ; n1996
g1355 and n1995_not n1996_not ; n1997
g1356 and n1994_not n1997 ; n1998
g1357 and n1994 n1997_not ; n1999
g1358 and in3[86] n1792 ; n2000
g1359 and in2[86] n1792_not ; n2001
g1360 and n2000_not n2001_not ; n2002
g1361 and in1[86] n1787 ; n2003
g1362 and in0[86] n1787_not ; n2004
g1363 and n2003_not n2004_not ; n2005
g1364 and n2002_not n2005 ; n2006
g1365 and n1999_not n2006_not ; n2007
g1366 and in1[85] n1787 ; n2008
g1367 and in0[85] n1787_not ; n2009
g1368 and n2008_not n2009_not ; n2010
g1369 and in3[85] n1792 ; n2011
g1370 and in2[85] n1792_not ; n2012
g1371 and n2011_not n2012_not ; n2013
g1372 and n2010 n2013_not ; n2014
g1373 and in1[84] n1787 ; n2015
g1374 and in0[84] n1787_not ; n2016
g1375 and n2015_not n2016_not ; n2017
g1376 and in3[84] n1792 ; n2018
g1377 and in2[84] n1792_not ; n2019
g1378 and n2018_not n2019_not ; n2020
g1379 and n2017_not n2020 ; n2021
g1380 and n2014_not n2021 ; n2022
g1381 and n2010_not n2013 ; n2023
g1382 and n2022_not n2023_not ; n2024
g1383 and n2007 n2024_not ; n2025
g1384 and n2002 n2005_not ; n2026
g1385 and n1999_not n2026 ; n2027
g1386 and in3[80] n1792 ; n2028
g1387 and in2[80] n1792_not ; n2029
g1388 and n2028_not n2029_not ; n2030
g1389 and in1[80] n1787 ; n2031
g1390 and in0[80] n1787_not ; n2032
g1391 and n2031_not n2032_not ; n2033
g1392 and n2030_not n2033 ; n2034
g1393 and in1[83] n1787 ; n2035
g1394 and in0[83] n1787_not ; n2036
g1395 and n2035_not n2036_not ; n2037
g1396 and in3[83] n1792 ; n2038
g1397 and in2[83] n1792_not ; n2039
g1398 and n2038_not n2039_not ; n2040
g1399 and n2037 n2040_not ; n2041
g1400 and in3[82] n1792 ; n2042
g1401 and in2[82] n1792_not ; n2043
g1402 and n2042_not n2043_not ; n2044
g1403 and in1[82] n1787 ; n2045
g1404 and in0[82] n1787_not ; n2046
g1405 and n2045_not n2046_not ; n2047
g1406 and n2044_not n2047 ; n2048
g1407 and n2041_not n2048_not ; n2049
g1408 and in1[81] n1787 ; n2050
g1409 and in0[81] n1787_not ; n2051
g1410 and n2050_not n2051_not ; n2052
g1411 and in3[81] n1792 ; n2053
g1412 and in2[81] n1792_not ; n2054
g1413 and n2053_not n2054_not ; n2055
g1414 and n2052 n2055_not ; n2056
g1415 and in1[79] n1787 ; n2057
g1416 and in0[79] n1787_not ; n2058
g1417 and n2057_not n2058_not ; n2059
g1418 and in3[79] n1792 ; n2060
g1419 and in2[79] n1792_not ; n2061
g1420 and n2060_not n2061_not ; n2062
g1421 and n2059_not n2062 ; n2063
g1422 and n2059 n2062_not ; n2064
g1423 and in3[78] n1792 ; n2065
g1424 and in2[78] n1792_not ; n2066
g1425 and n2065_not n2066_not ; n2067
g1426 and in1[78] n1787 ; n2068
g1427 and in0[78] n1787_not ; n2069
g1428 and n2068_not n2069_not ; n2070
g1429 and n2067_not n2070 ; n2071
g1430 and n2064_not n2071_not ; n2072
g1431 and in1[77] n1787 ; n2073
g1432 and in0[77] n1787_not ; n2074
g1433 and n2073_not n2074_not ; n2075
g1434 and in3[77] n1792 ; n2076
g1435 and in2[77] n1792_not ; n2077
g1436 and n2076_not n2077_not ; n2078
g1437 and n2075 n2078_not ; n2079
g1438 and in1[76] n1787 ; n2080
g1439 and in0[76] n1787_not ; n2081
g1440 and n2080_not n2081_not ; n2082
g1441 and in3[76] n1792 ; n2083
g1442 and in2[76] n1792_not ; n2084
g1443 and n2083_not n2084_not ; n2085
g1444 and n2082_not n2085 ; n2086
g1445 and n2079_not n2086 ; n2087
g1446 and n2075_not n2078 ; n2088
g1447 and n2087_not n2088_not ; n2089
g1448 and n2072 n2089_not ; n2090
g1449 and n2067 n2070_not ; n2091
g1450 and n2064_not n2091 ; n2092
g1451 and in1[71] n1787 ; n2093
g1452 and in0[71] n1787_not ; n2094
g1453 and n2093_not n2094_not ; n2095
g1454 and in3[71] n1792 ; n2096
g1455 and in2[71] n1792_not ; n2097
g1456 and n2096_not n2097_not ; n2098
g1457 and n2095_not n2098 ; n2099
g1458 and n2095 n2098_not ; n2100
g1459 and in3[70] n1792 ; n2101
g1460 and in2[70] n1792_not ; n2102
g1461 and n2101_not n2102_not ; n2103
g1462 and in1[70] n1787 ; n2104
g1463 and in0[70] n1787_not ; n2105
g1464 and n2104_not n2105_not ; n2106
g1465 and n2103_not n2106 ; n2107
g1466 and n2100_not n2107_not ; n2108
g1467 and in1[69] n1787 ; n2109
g1468 and in0[69] n1787_not ; n2110
g1469 and n2109_not n2110_not ; n2111
g1470 and in3[69] n1792 ; n2112
g1471 and in2[69] n1792_not ; n2113
g1472 and n2112_not n2113_not ; n2114
g1473 and n2111 n2114_not ; n2115
g1474 and in1[68] n1787 ; n2116
g1475 and in0[68] n1787_not ; n2117
g1476 and n2116_not n2117_not ; n2118
g1477 and in3[68] n1792 ; n2119
g1478 and in2[68] n1792_not ; n2120
g1479 and n2119_not n2120_not ; n2121
g1480 and n2118_not n2121 ; n2122
g1481 and n2115_not n2122 ; n2123
g1482 and n2111_not n2114 ; n2124
g1483 and n2123_not n2124_not ; n2125
g1484 and n2108 n2125_not ; n2126
g1485 and n2103 n2106_not ; n2127
g1486 and n2100_not n2127 ; n2128
g1487 and in1[67] n1787 ; n2129
g1488 and in0[67] n1787_not ; n2130
g1489 and n2129_not n2130_not ; n2131
g1490 and in3[67] n1792 ; n2132
g1491 and in2[67] n1792_not ; n2133
g1492 and n2132_not n2133_not ; n2134
g1493 and n2131 n2134_not ; n2135
g1494 and in3[66] n1792 ; n2136
g1495 and in2[66] n1792_not ; n2137
g1496 and n2136_not n2137_not ; n2138
g1497 and in1[66] n1787 ; n2139
g1498 and in0[66] n1787_not ; n2140
g1499 and n2139_not n2140_not ; n2141
g1500 and n2138_not n2141 ; n2142
g1501 and n2135_not n2142_not ; n2143
g1502 and in3[64] n1792 ; n2144
g1503 and in2[64] n1792_not ; n2145
g1504 and n2144_not n2145_not ; n2146
g1505 and in1[64] n1787 ; n2147
g1506 and in0[64] n1787_not ; n2148
g1507 and n2147_not n2148_not ; n2149
g1508 and n2146_not n2149 ; n2150
g1509 and in1[65] n1787 ; n2151
g1510 and in0[65] n1787_not ; n2152
g1511 and n2151_not n2152_not ; n2153
g1512 and in3[65] n1792 ; n2154
g1513 and in2[65] n1792_not ; n2155
g1514 and n2154_not n2155_not ; n2156
g1515 and n2153 n2156_not ; n2157
g1516 and in1[63] n1787 ; n2158
g1517 and in0[63] n1787_not ; n2159
g1518 and n2158_not n2159_not ; n2160
g1519 and in3[63] n1792 ; n2161
g1520 and in2[63] n1792_not ; n2162
g1521 and n2161_not n2162_not ; n2163
g1522 and n2160_not n2163 ; n2164
g1523 and n2160 n2163_not ; n2165
g1524 and in3[62] n1792 ; n2166
g1525 and in2[62] n1792_not ; n2167
g1526 and n2166_not n2167_not ; n2168
g1527 and in1[62] n1787 ; n2169
g1528 and in0[62] n1787_not ; n2170
g1529 and n2169_not n2170_not ; n2171
g1530 and n2168_not n2171 ; n2172
g1531 and n2165_not n2172_not ; n2173
g1532 and in1[60] n1787 ; n2174
g1533 and in0[60] n1787_not ; n2175
g1534 and n2174_not n2175_not ; n2176
g1535 and in3[60] n1792 ; n2177
g1536 and in2[60] n1792_not ; n2178
g1537 and n2177_not n2178_not ; n2179
g1538 and n2176 n2179_not ; n2180
g1539 and in1[61] n1787 ; n2181
g1540 and in0[61] n1787_not ; n2182
g1541 and n2181_not n2182_not ; n2183
g1542 and in3[61] n1792 ; n2184
g1543 and in2[61] n1792_not ; n2185
g1544 and n2184_not n2185_not ; n2186
g1545 and n2183 n2186_not ; n2187
g1546 and n2180_not n2187_not ; n2188
g1547 and n2173 n2188 ; n2189
g1548 and in1[59] n1787 ; n2190
g1549 and in0[59] n1787_not ; n2191
g1550 and n2190_not n2191_not ; n2192
g1551 and in3[59] n1792 ; n2193
g1552 and in2[59] n1792_not ; n2194
g1553 and n2193_not n2194_not ; n2195
g1554 and n2192_not n2195 ; n2196
g1555 and n2192 n2195_not ; n2197
g1556 and in1[58] n1787 ; n2198
g1557 and in0[58] n1787_not ; n2199
g1558 and n2198_not n2199_not ; n2200
g1559 and in3[58] n1792 ; n2201
g1560 and in2[58] n1792_not ; n2202
g1561 and n2201_not n2202_not ; n2203
g1562 and n2200 n2203_not ; n2204
g1563 and n2197_not n2204_not ; n2205
g1564 and in1[57] n1787 ; n2206
g1565 and in0[57] n1787_not ; n2207
g1566 and n2206_not n2207_not ; n2208
g1567 and in3[57] n1792 ; n2209
g1568 and in2[57] n1792_not ; n2210
g1569 and n2209_not n2210_not ; n2211
g1570 and n2208 n2211_not ; n2212
g1571 and in1[56] n1787 ; n2213
g1572 and in0[56] n1787_not ; n2214
g1573 and n2213_not n2214_not ; n2215
g1574 and in3[56] n1792 ; n2216
g1575 and in2[56] n1792_not ; n2217
g1576 and n2216_not n2217_not ; n2218
g1577 and n2215_not n2218 ; n2219
g1578 and n2212_not n2219 ; n2220
g1579 and n2208_not n2211 ; n2221
g1580 and n2220_not n2221_not ; n2222
g1581 and n2200_not n2203 ; n2223
g1582 and n2222 n2223_not ; n2224
g1583 and n2205 n2224_not ; n2225
g1584 and n2196_not n2225_not ; n2226
g1585 and n2189 n2226_not ; n2227
g1586 and n2176_not n2179 ; n2228
g1587 and n2187_not n2228 ; n2229
g1588 and n2183_not n2186 ; n2230
g1589 and n2229_not n2230_not ; n2231
g1590 and n2173 n2231_not ; n2232
g1591 and n2168 n2171_not ; n2233
g1592 and n2165_not n2233 ; n2234
g1593 and in1[47] n1787 ; n2235
g1594 and in0[47] n1787_not ; n2236
g1595 and n2235_not n2236_not ; n2237
g1596 and in3[47] n1792 ; n2238
g1597 and in2[47] n1792_not ; n2239
g1598 and n2238_not n2239_not ; n2240
g1599 and n2237_not n2240 ; n2241
g1600 and n2237 n2240_not ; n2242
g1601 and in3[46] n1792 ; n2243
g1602 and in2[46] n1792_not ; n2244
g1603 and n2243_not n2244_not ; n2245
g1604 and in1[46] n1787 ; n2246
g1605 and in0[46] n1787_not ; n2247
g1606 and n2246_not n2247_not ; n2248
g1607 and n2245_not n2248 ; n2249
g1608 and n2242_not n2249_not ; n2250
g1609 and in1[44] n1787 ; n2251
g1610 and in0[44] n1787_not ; n2252
g1611 and n2251_not n2252_not ; n2253
g1612 and in3[44] n1792 ; n2254
g1613 and in2[44] n1792_not ; n2255
g1614 and n2254_not n2255_not ; n2256
g1615 and n2253 n2256_not ; n2257
g1616 and in1[45] n1787 ; n2258
g1617 and in0[45] n1787_not ; n2259
g1618 and n2258_not n2259_not ; n2260
g1619 and in3[45] n1792 ; n2261
g1620 and in2[45] n1792_not ; n2262
g1621 and n2261_not n2262_not ; n2263
g1622 and n2260 n2263_not ; n2264
g1623 and n2257_not n2264_not ; n2265
g1624 and n2250 n2265 ; n2266
g1625 and in1[43] n1787 ; n2267
g1626 and in0[43] n1787_not ; n2268
g1627 and n2267_not n2268_not ; n2269
g1628 and in3[43] n1792 ; n2270
g1629 and in2[43] n1792_not ; n2271
g1630 and n2270_not n2271_not ; n2272
g1631 and n2269_not n2272 ; n2273
g1632 and n2269 n2272_not ; n2274
g1633 and in1[42] n1787 ; n2275
g1634 and in0[42] n1787_not ; n2276
g1635 and n2275_not n2276_not ; n2277
g1636 and in3[42] n1792 ; n2278
g1637 and in2[42] n1792_not ; n2279
g1638 and n2278_not n2279_not ; n2280
g1639 and n2277 n2280_not ; n2281
g1640 and n2274_not n2281_not ; n2282
g1641 and in1[41] n1787 ; n2283
g1642 and in0[41] n1787_not ; n2284
g1643 and n2283_not n2284_not ; n2285
g1644 and in3[41] n1792 ; n2286
g1645 and in2[41] n1792_not ; n2287
g1646 and n2286_not n2287_not ; n2288
g1647 and n2285 n2288_not ; n2289
g1648 and in1[40] n1787 ; n2290
g1649 and in0[40] n1787_not ; n2291
g1650 and n2290_not n2291_not ; n2292
g1651 and in3[40] n1792 ; n2293
g1652 and in2[40] n1792_not ; n2294
g1653 and n2293_not n2294_not ; n2295
g1654 and n2292_not n2295 ; n2296
g1655 and n2289_not n2296 ; n2297
g1656 and n2285_not n2288 ; n2298
g1657 and n2297_not n2298_not ; n2299
g1658 and n2277_not n2280 ; n2300
g1659 and n2299 n2300_not ; n2301
g1660 and n2282 n2301_not ; n2302
g1661 and n2273_not n2302_not ; n2303
g1662 and n2266 n2303_not ; n2304
g1663 and n2253_not n2256 ; n2305
g1664 and n2264_not n2305 ; n2306
g1665 and n2260_not n2263 ; n2307
g1666 and n2306_not n2307_not ; n2308
g1667 and n2250 n2308_not ; n2309
g1668 and n2245 n2248_not ; n2310
g1669 and n2242_not n2310 ; n2311
g1670 and in3[32] n1792 ; n2312
g1671 and in2[32] n1792_not ; n2313
g1672 and n2312_not n2313_not ; n2314
g1673 and in1[32] n1787 ; n2315
g1674 and in0[32] n1787_not ; n2316
g1675 and n2315_not n2316_not ; n2317
g1676 and n2314_not n2317 ; n2318
g1677 and in1[31] n1787 ; n2319
g1678 and in0[31] n1787_not ; n2320
g1679 and n2319_not n2320_not ; n2321
g1680 and in3[31] n1792 ; n2322
g1681 and in2[31] n1792_not ; n2323
g1682 and n2322_not n2323_not ; n2324
g1683 and n2321 n2324_not ; n2325
g1684 and in1[30] n1787 ; n2326
g1685 and in0[30] n1787_not ; n2327
g1686 and n2326_not n2327_not ; n2328
g1687 and in3[30] n1792 ; n2329
g1688 and in2[30] n1792_not ; n2330
g1689 and n2329_not n2330_not ; n2331
g1690 and n2328 n2331_not ; n2332
g1691 and in1[29] n1787 ; n2333
g1692 and in0[29] n1787_not ; n2334
g1693 and n2333_not n2334_not ; n2335
g1694 and in3[29] n1792 ; n2336
g1695 and in2[29] n1792_not ; n2337
g1696 and n2336_not n2337_not ; n2338
g1697 and n2335 n2338_not ; n2339
g1698 and in1[28] n1787 ; n2340
g1699 and in0[28] n1787_not ; n2341
g1700 and n2340_not n2341_not ; n2342
g1701 and in3[28] n1792 ; n2343
g1702 and in2[28] n1792_not ; n2344
g1703 and n2343_not n2344_not ; n2345
g1704 and n2342 n2345_not ; n2346
g1705 and in1[27] n1787 ; n2347
g1706 and in0[27] n1787_not ; n2348
g1707 and n2347_not n2348_not ; n2349
g1708 and in3[27] n1792 ; n2350
g1709 and in2[27] n1792_not ; n2351
g1710 and n2350_not n2351_not ; n2352
g1711 and n2349 n2352_not ; n2353
g1712 and in1[26] n1787 ; n2354
g1713 and in0[26] n1787_not ; n2355
g1714 and n2354_not n2355_not ; n2356
g1715 and in3[26] n1792 ; n2357
g1716 and in2[26] n1792_not ; n2358
g1717 and n2357_not n2358_not ; n2359
g1718 and n2356 n2359_not ; n2360
g1719 and in3[25] n1792 ; n2361
g1720 and in2[25] n1792_not ; n2362
g1721 and n2361_not n2362_not ; n2363
g1722 and in3[24] n1792 ; n2364
g1723 and in2[24] n1792_not ; n2365
g1724 and n2364_not n2365_not ; n2366
g1725 and in1[23] n1787 ; n2367
g1726 and in0[23] n1787_not ; n2368
g1727 and n2367_not n2368_not ; n2369
g1728 and in3[23] n1792 ; n2370
g1729 and in2[23] n1792_not ; n2371
g1730 and n2370_not n2371_not ; n2372
g1731 and n2369 n2372_not ; n2373
g1732 and in1[22] n1787 ; n2374
g1733 and in0[22] n1787_not ; n2375
g1734 and n2374_not n2375_not ; n2376
g1735 and in3[22] n1792 ; n2377
g1736 and in2[22] n1792_not ; n2378
g1737 and n2377_not n2378_not ; n2379
g1738 and n2376 n2379_not ; n2380
g1739 and in1[21] n1787 ; n2381
g1740 and in0[21] n1787_not ; n2382
g1741 and n2381_not n2382_not ; n2383
g1742 and in3[21] n1792 ; n2384
g1743 and in2[21] n1792_not ; n2385
g1744 and n2384_not n2385_not ; n2386
g1745 and n2383 n2386_not ; n2387
g1746 and in1[20] n1787 ; n2388
g1747 and in0[20] n1787_not ; n2389
g1748 and n2388_not n2389_not ; n2390
g1749 and in3[20] n1792 ; n2391
g1750 and in2[20] n1792_not ; n2392
g1751 and n2391_not n2392_not ; n2393
g1752 and n2390 n2393_not ; n2394
g1753 and in1[19] n1787 ; n2395
g1754 and in0[19] n1787_not ; n2396
g1755 and n2395_not n2396_not ; n2397
g1756 and in3[19] n1792 ; n2398
g1757 and in2[19] n1792_not ; n2399
g1758 and n2398_not n2399_not ; n2400
g1759 and n2397 n2400_not ; n2401
g1760 and in1[18] n1787 ; n2402
g1761 and in0[18] n1787_not ; n2403
g1762 and n2402_not n2403_not ; n2404
g1763 and in3[18] n1792 ; n2405
g1764 and in2[18] n1792_not ; n2406
g1765 and n2405_not n2406_not ; n2407
g1766 and n2404 n2407_not ; n2408
g1767 and in3[17] n1792 ; n2409
g1768 and in2[17] n1792_not ; n2410
g1769 and n2409_not n2410_not ; n2411
g1770 and in3[16] n1792 ; n2412
g1771 and in2[16] n1792_not ; n2413
g1772 and n2412_not n2413_not ; n2414
g1773 and in1[15] n1787 ; n2415
g1774 and in0[15] n1787_not ; n2416
g1775 and n2415_not n2416_not ; n2417
g1776 and in3[15] n1792 ; n2418
g1777 and in2[15] n1792_not ; n2419
g1778 and n2418_not n2419_not ; n2420
g1779 and n2417 n2420_not ; n2421
g1780 and in1[14] n1787 ; n2422
g1781 and in0[14] n1787_not ; n2423
g1782 and n2422_not n2423_not ; n2424
g1783 and in3[14] n1792 ; n2425
g1784 and in2[14] n1792_not ; n2426
g1785 and n2425_not n2426_not ; n2427
g1786 and n2424 n2427_not ; n2428
g1787 and in1[13] n1787 ; n2429
g1788 and in0[13] n1787_not ; n2430
g1789 and n2429_not n2430_not ; n2431
g1790 and in3[13] n1792 ; n2432
g1791 and in2[13] n1792_not ; n2433
g1792 and n2432_not n2433_not ; n2434
g1793 and n2431 n2434_not ; n2435
g1794 and in1[12] n1787 ; n2436
g1795 and in0[12] n1787_not ; n2437
g1796 and n2436_not n2437_not ; n2438
g1797 and in3[12] n1792 ; n2439
g1798 and in2[12] n1792_not ; n2440
g1799 and n2439_not n2440_not ; n2441
g1800 and n2438 n2441_not ; n2442
g1801 and in1[11] n1787 ; n2443
g1802 and in0[11] n1787_not ; n2444
g1803 and n2443_not n2444_not ; n2445
g1804 and in3[11] n1792 ; n2446
g1805 and in2[11] n1792_not ; n2447
g1806 and n2446_not n2447_not ; n2448
g1807 and n2445 n2448_not ; n2449
g1808 and in1[10] n1787 ; n2450
g1809 and in0[10] n1787_not ; n2451
g1810 and n2450_not n2451_not ; n2452
g1811 and in3[10] n1792 ; n2453
g1812 and in2[10] n1792_not ; n2454
g1813 and n2453_not n2454_not ; n2455
g1814 and n2452 n2455_not ; n2456
g1815 and in3[9] n1792 ; n2457
g1816 and in2[9] n1792_not ; n2458
g1817 and n2457_not n2458_not ; n2459
g1818 and in3[8] n1792 ; n2460
g1819 and in2[8] n1792_not ; n2461
g1820 and n2460_not n2461_not ; n2462
g1821 and in1[7] n1787 ; n2463
g1822 and in0[7] n1787_not ; n2464
g1823 and n2463_not n2464_not ; n2465
g1824 and in3[7] n1792 ; n2466
g1825 and in2[7] n1792_not ; n2467
g1826 and n2466_not n2467_not ; n2468
g1827 and n2465 n2468_not ; n2469
g1828 and in3[6] n1792 ; n2470
g1829 and in2[6] n1792_not ; n2471
g1830 and n2470_not n2471_not ; n2472
g1831 and in1[6] n1787 ; n2473
g1832 and in0[6] n1787_not ; n2474
g1833 and n2473_not n2474_not ; n2475
g1834 and in3[5] n1792 ; n2476
g1835 and in2[5] n1792_not ; n2477
g1836 and n2476_not n2477_not ; n2478
g1837 and in1[5] n1787 ; n2479
g1838 and in0[5] n1787_not ; n2480
g1839 and n2479_not n2480_not ; n2481
g1840 and in3[4] n1792 ; n2482
g1841 and in2[4] n1792_not ; n2483
g1842 and n2482_not n2483_not ; n2484
g1843 and in1[4] n1787 ; n2485
g1844 and in0[4] n1787_not ; n2486
g1845 and n2485_not n2486_not ; n2487
g1846 and in1[3] n1787 ; n2488
g1847 and in0[3] n1787_not ; n2489
g1848 and n2488_not n2489_not ; n2490
g1849 and in3[3] n1792 ; n2491
g1850 and in2[3] n1792_not ; n2492
g1851 and n2491_not n2492_not ; n2493
g1852 and n2490 n2493_not ; n2494
g1853 and in3[1] n1792 ; n2495
g1854 and in2[1] n1792_not ; n2496
g1855 and n2495_not n2496_not ; n2497
g1856 and in1[0] n1787 ; n2498
g1857 and in0[0] n1787_not ; n2499
g1858 and n2498_not n2499_not ; n2500
g1859 and in3[0] n1792 ; n2501
g1860 and in2[0] n1792_not ; n2502
g1861 and n2501_not n2502_not ; n2503
g1862 and n2500_not n2503 ; n2504
g1863 and n2497 n2504 ; n2505
g1864 and in1[1] n1787 ; n2506
g1865 and in0[1] n1787_not ; n2507
g1866 and n2506_not n2507_not ; n2508
g1867 and n2505_not n2508 ; n2509
g1868 and in1[2] n1787 ; n2510
g1869 and in0[2] n1787_not ; n2511
g1870 and n2510_not n2511_not ; n2512
g1871 and in3[2] n1792 ; n2513
g1872 and in2[2] n1792_not ; n2514
g1873 and n2513_not n2514_not ; n2515
g1874 and n2512 n2515_not ; n2516
g1875 and n2497_not n2504_not ; n2517
g1876 and n2516_not n2517_not ; n2518
g1877 and n2509_not n2518 ; n2519
g1878 and n2512_not n2515 ; n2520
g1879 and n2519_not n2520_not ; n2521
g1880 and n2494_not n2521_not ; n2522
g1881 and n2490_not n2493 ; n2523
g1882 and n2522_not n2523_not ; n2524
g1883 and n2487 n2524 ; n2525
g1884 and n2484 n2525_not ; n2526
g1885 and n2487_not n2524_not ; n2527
g1886 and n2526_not n2527_not ; n2528
g1887 and n2481 n2528 ; n2529
g1888 and n2478 n2529_not ; n2530
g1889 and n2481_not n2528_not ; n2531
g1890 and n2530_not n2531_not ; n2532
g1891 and n2475 n2532 ; n2533
g1892 and n2472 n2533_not ; n2534
g1893 and n2475_not n2532_not ; n2535
g1894 and n2534_not n2535_not ; n2536
g1895 and n2469_not n2536_not ; n2537
g1896 and n2465_not n2468 ; n2538
g1897 and n2537_not n2538_not ; n2539
g1898 and in1[8] n1787 ; n2540
g1899 and in0[8] n1787_not ; n2541
g1900 and n2540_not n2541_not ; n2542
g1901 and n2539 n2542 ; n2543
g1902 and n2462 n2543_not ; n2544
g1903 and n2539_not n2542_not ; n2545
g1904 and n2544_not n2545_not ; n2546
g1905 and in1[9] n1787 ; n2547
g1906 and in0[9] n1787_not ; n2548
g1907 and n2547_not n2548_not ; n2549
g1908 and n2546 n2549 ; n2550
g1909 and n2459 n2550_not ; n2551
g1910 and n2546_not n2549_not ; n2552
g1911 and n2551_not n2552_not ; n2553
g1912 and n2456_not n2553_not ; n2554
g1913 and n2452_not n2455 ; n2555
g1914 and n2554_not n2555_not ; n2556
g1915 and n2449_not n2556_not ; n2557
g1916 and n2445_not n2448 ; n2558
g1917 and n2557_not n2558_not ; n2559
g1918 and n2442_not n2559_not ; n2560
g1919 and n2438_not n2441 ; n2561
g1920 and n2560_not n2561_not ; n2562
g1921 and n2435_not n2562_not ; n2563
g1922 and n2431_not n2434 ; n2564
g1923 and n2563_not n2564_not ; n2565
g1924 and n2428_not n2565_not ; n2566
g1925 and n2424_not n2427 ; n2567
g1926 and n2566_not n2567_not ; n2568
g1927 and n2421_not n2568_not ; n2569
g1928 and n2417_not n2420 ; n2570
g1929 and n2569_not n2570_not ; n2571
g1930 and in1[16] n1787 ; n2572
g1931 and in0[16] n1787_not ; n2573
g1932 and n2572_not n2573_not ; n2574
g1933 and n2571 n2574 ; n2575
g1934 and n2414 n2575_not ; n2576
g1935 and n2571_not n2574_not ; n2577
g1936 and n2576_not n2577_not ; n2578
g1937 and in1[17] n1787 ; n2579
g1938 and in0[17] n1787_not ; n2580
g1939 and n2579_not n2580_not ; n2581
g1940 and n2578 n2581 ; n2582
g1941 and n2411 n2582_not ; n2583
g1942 and n2578_not n2581_not ; n2584
g1943 and n2583_not n2584_not ; n2585
g1944 and n2408_not n2585_not ; n2586
g1945 and n2404_not n2407 ; n2587
g1946 and n2586_not n2587_not ; n2588
g1947 and n2401_not n2588_not ; n2589
g1948 and n2397_not n2400 ; n2590
g1949 and n2589_not n2590_not ; n2591
g1950 and n2394_not n2591_not ; n2592
g1951 and n2390_not n2393 ; n2593
g1952 and n2592_not n2593_not ; n2594
g1953 and n2387_not n2594_not ; n2595
g1954 and n2383_not n2386 ; n2596
g1955 and n2595_not n2596_not ; n2597
g1956 and n2380_not n2597_not ; n2598
g1957 and n2376_not n2379 ; n2599
g1958 and n2598_not n2599_not ; n2600
g1959 and n2373_not n2600_not ; n2601
g1960 and n2369_not n2372 ; n2602
g1961 and n2601_not n2602_not ; n2603
g1962 and in1[24] n1787 ; n2604
g1963 and in0[24] n1787_not ; n2605
g1964 and n2604_not n2605_not ; n2606
g1965 and n2603 n2606 ; n2607
g1966 and n2366 n2607_not ; n2608
g1967 and n2603_not n2606_not ; n2609
g1968 and n2608_not n2609_not ; n2610
g1969 and in1[25] n1787 ; n2611
g1970 and in0[25] n1787_not ; n2612
g1971 and n2611_not n2612_not ; n2613
g1972 and n2610 n2613 ; n2614
g1973 and n2363 n2614_not ; n2615
g1974 and n2610_not n2613_not ; n2616
g1975 and n2615_not n2616_not ; n2617
g1976 and n2360_not n2617_not ; n2618
g1977 and n2356_not n2359 ; n2619
g1978 and n2618_not n2619_not ; n2620
g1979 and n2353_not n2620_not ; n2621
g1980 and n2349_not n2352 ; n2622
g1981 and n2621_not n2622_not ; n2623
g1982 and n2346_not n2623_not ; n2624
g1983 and n2342_not n2345 ; n2625
g1984 and n2624_not n2625_not ; n2626
g1985 and n2339_not n2626_not ; n2627
g1986 and n2335_not n2338 ; n2628
g1987 and n2627_not n2628_not ; n2629
g1988 and n2332_not n2629_not ; n2630
g1989 and n2328_not n2331 ; n2631
g1990 and n2630_not n2631_not ; n2632
g1991 and n2325_not n2632_not ; n2633
g1992 and n2321_not n2324 ; n2634
g1993 and n2633_not n2634_not ; n2635
g1994 and in1[39] n1787 ; n2636
g1995 and in0[39] n1787_not ; n2637
g1996 and n2636_not n2637_not ; n2638
g1997 and in3[39] n1792 ; n2639
g1998 and in2[39] n1792_not ; n2640
g1999 and n2639_not n2640_not ; n2641
g2000 and n2638 n2641_not ; n2642
g2001 and in3[38] n1792 ; n2643
g2002 and in2[38] n1792_not ; n2644
g2003 and n2643_not n2644_not ; n2645
g2004 and in1[38] n1787 ; n2646
g2005 and in0[38] n1787_not ; n2647
g2006 and n2646_not n2647_not ; n2648
g2007 and n2645_not n2648 ; n2649
g2008 and n2642_not n2649_not ; n2650
g2009 and in1[36] n1787 ; n2651
g2010 and in0[36] n1787_not ; n2652
g2011 and n2651_not n2652_not ; n2653
g2012 and in3[36] n1792 ; n2654
g2013 and in2[36] n1792_not ; n2655
g2014 and n2654_not n2655_not ; n2656
g2015 and n2653 n2656_not ; n2657
g2016 and in1[37] n1787 ; n2658
g2017 and in0[37] n1787_not ; n2659
g2018 and n2658_not n2659_not ; n2660
g2019 and in3[37] n1792 ; n2661
g2020 and in2[37] n1792_not ; n2662
g2021 and n2661_not n2662_not ; n2663
g2022 and n2660 n2663_not ; n2664
g2023 and n2657_not n2664_not ; n2665
g2024 and n2650 n2665 ; n2666
g2025 and in1[33] n1787 ; n2667
g2026 and in0[33] n1787_not ; n2668
g2027 and n2667_not n2668_not ; n2669
g2028 and in3[33] n1792 ; n2670
g2029 and in2[33] n1792_not ; n2671
g2030 and n2670_not n2671_not ; n2672
g2031 and n2669 n2672_not ; n2673
g2032 and in1[35] n1787 ; n2674
g2033 and in0[35] n1787_not ; n2675
g2034 and n2674_not n2675_not ; n2676
g2035 and in3[35] n1792 ; n2677
g2036 and in2[35] n1792_not ; n2678
g2037 and n2677_not n2678_not ; n2679
g2038 and n2676 n2679_not ; n2680
g2039 and in3[34] n1792 ; n2681
g2040 and in2[34] n1792_not ; n2682
g2041 and n2681_not n2682_not ; n2683
g2042 and in1[34] n1787 ; n2684
g2043 and in0[34] n1787_not ; n2685
g2044 and n2684_not n2685_not ; n2686
g2045 and n2683_not n2686 ; n2687
g2046 and n2680_not n2687_not ; n2688
g2047 and n2673_not n2688 ; n2689
g2048 and n2666 n2689 ; n2690
g2049 and n2635_not n2690 ; n2691
g2050 and n2318_not n2691 ; n2692
g2051 and n2638_not n2641 ; n2693
g2052 and n2653_not n2656 ; n2694
g2053 and n2664_not n2694 ; n2695
g2054 and n2660_not n2663 ; n2696
g2055 and n2695_not n2696_not ; n2697
g2056 and n2650 n2697_not ; n2698
g2057 and n2642_not n2645 ; n2699
g2058 and n2648_not n2699 ; n2700
g2059 and n2676_not n2679 ; n2701
g2060 and n2680_not n2683 ; n2702
g2061 and n2686_not n2702 ; n2703
g2062 and n2314 n2317_not ; n2704
g2063 and n2669_not n2672 ; n2705
g2064 and n2704_not n2705_not ; n2706
g2065 and n2689 n2706_not ; n2707
g2066 and n2703_not n2707_not ; n2708
g2067 and n2701_not n2708 ; n2709
g2068 and n2666 n2709_not ; n2710
g2069 and n2700_not n2710_not ; n2711
g2070 and n2698_not n2711 ; n2712
g2071 and n2693_not n2712 ; n2713
g2072 and n2692_not n2713 ; n2714
g2073 and n2292 n2295_not ; n2715
g2074 and n2289_not n2715_not ; n2716
g2075 and n2282 n2716 ; n2717
g2076 and n2266 n2717 ; n2718
g2077 and n2714_not n2718 ; n2719
g2078 and n2311_not n2719_not ; n2720
g2079 and n2309_not n2720 ; n2721
g2080 and n2304_not n2721 ; n2722
g2081 and n2241_not n2722 ; n2723
g2082 and in3[48] n1792 ; n2724
g2083 and in2[48] n1792_not ; n2725
g2084 and n2724_not n2725_not ; n2726
g2085 and in1[48] n1787 ; n2727
g2086 and in0[48] n1787_not ; n2728
g2087 and n2727_not n2728_not ; n2729
g2088 and n2726_not n2729 ; n2730
g2089 and in1[55] n1787 ; n2731
g2090 and in0[55] n1787_not ; n2732
g2091 and n2731_not n2732_not ; n2733
g2092 and in3[55] n1792 ; n2734
g2093 and in2[55] n1792_not ; n2735
g2094 and n2734_not n2735_not ; n2736
g2095 and n2733 n2736_not ; n2737
g2096 and in3[54] n1792 ; n2738
g2097 and in2[54] n1792_not ; n2739
g2098 and n2738_not n2739_not ; n2740
g2099 and in1[54] n1787 ; n2741
g2100 and in0[54] n1787_not ; n2742
g2101 and n2741_not n2742_not ; n2743
g2102 and n2740_not n2743 ; n2744
g2103 and n2737_not n2744_not ; n2745
g2104 and in1[53] n1787 ; n2746
g2105 and in0[53] n1787_not ; n2747
g2106 and n2746_not n2747_not ; n2748
g2107 and in3[53] n1792 ; n2749
g2108 and in2[53] n1792_not ; n2750
g2109 and n2749_not n2750_not ; n2751
g2110 and n2748 n2751_not ; n2752
g2111 and in3[52] n1792 ; n2753
g2112 and in2[52] n1792_not ; n2754
g2113 and n2753_not n2754_not ; n2755
g2114 and in1[52] n1787 ; n2756
g2115 and in0[52] n1787_not ; n2757
g2116 and n2756_not n2757_not ; n2758
g2117 and n2755_not n2758 ; n2759
g2118 and n2752_not n2759_not ; n2760
g2119 and n2745 n2760 ; n2761
g2120 and in1[49] n1787 ; n2762
g2121 and in0[49] n1787_not ; n2763
g2122 and n2762_not n2763_not ; n2764
g2123 and in3[49] n1792 ; n2765
g2124 and in2[49] n1792_not ; n2766
g2125 and n2765_not n2766_not ; n2767
g2126 and n2764 n2767_not ; n2768
g2127 and in1[51] n1787 ; n2769
g2128 and in0[51] n1787_not ; n2770
g2129 and n2769_not n2770_not ; n2771
g2130 and in3[51] n1792 ; n2772
g2131 and in2[51] n1792_not ; n2773
g2132 and n2772_not n2773_not ; n2774
g2133 and n2771 n2774_not ; n2775
g2134 and in3[50] n1792 ; n2776
g2135 and in2[50] n1792_not ; n2777
g2136 and n2776_not n2777_not ; n2778
g2137 and in1[50] n1787 ; n2779
g2138 and in0[50] n1787_not ; n2780
g2139 and n2779_not n2780_not ; n2781
g2140 and n2778_not n2781 ; n2782
g2141 and n2775_not n2782_not ; n2783
g2142 and n2768_not n2783 ; n2784
g2143 and n2761 n2784 ; n2785
g2144 and n2730_not n2785 ; n2786
g2145 and n2723_not n2786 ; n2787
g2146 and n2733_not n2736 ; n2788
g2147 and n2771_not n2774 ; n2789
g2148 and n2775_not n2778 ; n2790
g2149 and n2781_not n2790 ; n2791
g2150 and n2726 n2729_not ; n2792
g2151 and n2764_not n2767 ; n2793
g2152 and n2792_not n2793_not ; n2794
g2153 and n2784 n2794_not ; n2795
g2154 and n2791_not n2795_not ; n2796
g2155 and n2789_not n2796 ; n2797
g2156 and n2761 n2797_not ; n2798
g2157 and n2755 n2758_not ; n2799
g2158 and n2752_not n2799 ; n2800
g2159 and n2748_not n2751 ; n2801
g2160 and n2800_not n2801_not ; n2802
g2161 and n2740 n2743_not ; n2803
g2162 and n2802 n2803_not ; n2804
g2163 and n2745 n2804_not ; n2805
g2164 and n2798_not n2805_not ; n2806
g2165 and n2788_not n2806 ; n2807
g2166 and n2787_not n2807 ; n2808
g2167 and n2215 n2218_not ; n2809
g2168 and n2212_not n2809_not ; n2810
g2169 and n2189 n2810 ; n2811
g2170 and n2205 n2811 ; n2812
g2171 and n2808_not n2812 ; n2813
g2172 and n2234_not n2813_not ; n2814
g2173 and n2232_not n2814 ; n2815
g2174 and n2227_not n2815 ; n2816
g2175 and n2164_not n2816 ; n2817
g2176 and n2157_not n2817_not ; n2818
g2177 and n2150_not n2818 ; n2819
g2178 and n2143 n2819 ; n2820
g2179 and n2131_not n2134 ; n2821
g2180 and n2146 n2157_not ; n2822
g2181 and n2149_not n2822 ; n2823
g2182 and n2153_not n2156 ; n2824
g2183 and n2823_not n2824_not ; n2825
g2184 and n2138 n2141_not ; n2826
g2185 and n2825 n2826_not ; n2827
g2186 and n2143 n2827_not ; n2828
g2187 and n2821_not n2828_not ; n2829
g2188 and n2820_not n2829 ; n2830
g2189 and n2118 n2121_not ; n2831
g2190 and n2115_not n2831_not ; n2832
g2191 and n2108 n2832 ; n2833
g2192 and n2830_not n2833 ; n2834
g2193 and n2128_not n2834_not ; n2835
g2194 and n2126_not n2835 ; n2836
g2195 and n2099_not n2836 ; n2837
g2196 and in1[75] n1787 ; n2838
g2197 and in0[75] n1787_not ; n2839
g2198 and n2838_not n2839_not ; n2840
g2199 and in3[75] n1792 ; n2841
g2200 and in2[75] n1792_not ; n2842
g2201 and n2841_not n2842_not ; n2843
g2202 and n2840 n2843_not ; n2844
g2203 and in3[74] n1792 ; n2845
g2204 and in2[74] n1792_not ; n2846
g2205 and n2845_not n2846_not ; n2847
g2206 and in1[74] n1787 ; n2848
g2207 and in0[74] n1787_not ; n2849
g2208 and n2848_not n2849_not ; n2850
g2209 and n2847_not n2850 ; n2851
g2210 and n2844_not n2851_not ; n2852
g2211 and in1[73] n1787 ; n2853
g2212 and in0[73] n1787_not ; n2854
g2213 and n2853_not n2854_not ; n2855
g2214 and in3[73] n1792 ; n2856
g2215 and in2[73] n1792_not ; n2857
g2216 and n2856_not n2857_not ; n2858
g2217 and n2855 n2858_not ; n2859
g2218 and in3[72] n1792 ; n2860
g2219 and in2[72] n1792_not ; n2861
g2220 and n2860_not n2861_not ; n2862
g2221 and in1[72] n1787 ; n2863
g2222 and in0[72] n1787_not ; n2864
g2223 and n2863_not n2864_not ; n2865
g2224 and n2862_not n2865 ; n2866
g2225 and n2859_not n2866_not ; n2867
g2226 and n2852 n2867 ; n2868
g2227 and n2837_not n2868 ; n2869
g2228 and n2840_not n2843 ; n2870
g2229 and n2862 n2865_not ; n2871
g2230 and n2859_not n2871 ; n2872
g2231 and n2855_not n2858 ; n2873
g2232 and n2872_not n2873_not ; n2874
g2233 and n2847 n2850_not ; n2875
g2234 and n2874 n2875_not ; n2876
g2235 and n2852 n2876_not ; n2877
g2236 and n2870_not n2877_not ; n2878
g2237 and n2869_not n2878 ; n2879
g2238 and n2082 n2085_not ; n2880
g2239 and n2079_not n2880_not ; n2881
g2240 and n2072 n2881 ; n2882
g2241 and n2879_not n2882 ; n2883
g2242 and n2092_not n2883_not ; n2884
g2243 and n2090_not n2884 ; n2885
g2244 and n2063_not n2885 ; n2886
g2245 and n2056_not n2886_not ; n2887
g2246 and n2049 n2887 ; n2888
g2247 and n2034_not n2888 ; n2889
g2248 and n2037_not n2040 ; n2890
g2249 and n2030 n2056_not ; n2891
g2250 and n2033_not n2891 ; n2892
g2251 and n2052_not n2055 ; n2893
g2252 and n2892_not n2893_not ; n2894
g2253 and n2044 n2047_not ; n2895
g2254 and n2894 n2895_not ; n2896
g2255 and n2049 n2896_not ; n2897
g2256 and n2890_not n2897_not ; n2898
g2257 and n2889_not n2898 ; n2899
g2258 and n2017 n2020_not ; n2900
g2259 and n2014_not n2900_not ; n2901
g2260 and n2007 n2901 ; n2902
g2261 and n2899_not n2902 ; n2903
g2262 and n2027_not n2903_not ; n2904
g2263 and n2025_not n2904 ; n2905
g2264 and n1998_not n2905 ; n2906
g2265 and in1[91] n1787 ; n2907
g2266 and in0[91] n1787_not ; n2908
g2267 and n2907_not n2908_not ; n2909
g2268 and in3[91] n1792 ; n2910
g2269 and in2[91] n1792_not ; n2911
g2270 and n2910_not n2911_not ; n2912
g2271 and n2909 n2912_not ; n2913
g2272 and in3[90] n1792 ; n2914
g2273 and in2[90] n1792_not ; n2915
g2274 and n2914_not n2915_not ; n2916
g2275 and in1[90] n1787 ; n2917
g2276 and in0[90] n1787_not ; n2918
g2277 and n2917_not n2918_not ; n2919
g2278 and n2916_not n2919 ; n2920
g2279 and n2913_not n2920_not ; n2921
g2280 and in1[89] n1787 ; n2922
g2281 and in0[89] n1787_not ; n2923
g2282 and n2922_not n2923_not ; n2924
g2283 and in3[89] n1792 ; n2925
g2284 and in2[89] n1792_not ; n2926
g2285 and n2925_not n2926_not ; n2927
g2286 and n2924 n2927_not ; n2928
g2287 and in3[88] n1792 ; n2929
g2288 and in2[88] n1792_not ; n2930
g2289 and n2929_not n2930_not ; n2931
g2290 and in1[88] n1787 ; n2932
g2291 and in0[88] n1787_not ; n2933
g2292 and n2932_not n2933_not ; n2934
g2293 and n2931_not n2934 ; n2935
g2294 and n2928_not n2935_not ; n2936
g2295 and n2921 n2936 ; n2937
g2296 and n2906_not n2937 ; n2938
g2297 and n2909_not n2912 ; n2939
g2298 and n2931 n2934_not ; n2940
g2299 and n2928_not n2940 ; n2941
g2300 and n2924_not n2927 ; n2942
g2301 and n2941_not n2942_not ; n2943
g2302 and n2916 n2919_not ; n2944
g2303 and n2943 n2944_not ; n2945
g2304 and n2921 n2945_not ; n2946
g2305 and n2939_not n2946_not ; n2947
g2306 and n2938_not n2947 ; n2948
g2307 and n1981 n1984_not ; n2949
g2308 and n1978_not n2949_not ; n2950
g2309 and n1971 n2950 ; n2951
g2310 and n2948_not n2951 ; n2952
g2311 and n1991_not n2952_not ; n2953
g2312 and n1989_not n2953 ; n2954
g2313 and n1962_not n2954 ; n2955
g2314 and n1955_not n2955_not ; n2956
g2315 and n1948 n2956 ; n2957
g2316 and n1933_not n2957 ; n2958
g2317 and n1936_not n1939 ; n2959
g2318 and n1929 n1955_not ; n2960
g2319 and n1932_not n2960 ; n2961
g2320 and n1951_not n1954 ; n2962
g2321 and n2961_not n2962_not ; n2963
g2322 and n1943 n1946_not ; n2964
g2323 and n2963 n2964_not ; n2965
g2324 and n1948 n2965_not ; n2966
g2325 and n2959_not n2966_not ; n2967
g2326 and n2958_not n2967 ; n2968
g2327 and n1916 n1919_not ; n2969
g2328 and n1913_not n2969_not ; n2970
g2329 and n1906 n2970 ; n2971
g2330 and n2968_not n2971 ; n2972
g2331 and n1926_not n2972_not ; n2973
g2332 and n1924_not n2973 ; n2974
g2333 and n1897_not n2974 ; n2975
g2334 and in1[107] n1787 ; n2976
g2335 and in0[107] n1787_not ; n2977
g2336 and n2976_not n2977_not ; n2978
g2337 and in3[107] n1792 ; n2979
g2338 and in2[107] n1792_not ; n2980
g2339 and n2979_not n2980_not ; n2981
g2340 and n2978 n2981_not ; n2982
g2341 and in3[106] n1792 ; n2983
g2342 and in2[106] n1792_not ; n2984
g2343 and n2983_not n2984_not ; n2985
g2344 and in1[106] n1787 ; n2986
g2345 and in0[106] n1787_not ; n2987
g2346 and n2986_not n2987_not ; n2988
g2347 and n2985_not n2988 ; n2989
g2348 and n2982_not n2989_not ; n2990
g2349 and in1[105] n1787 ; n2991
g2350 and in0[105] n1787_not ; n2992
g2351 and n2991_not n2992_not ; n2993
g2352 and in3[105] n1792 ; n2994
g2353 and in2[105] n1792_not ; n2995
g2354 and n2994_not n2995_not ; n2996
g2355 and n2993 n2996_not ; n2997
g2356 and in3[104] n1792 ; n2998
g2357 and in2[104] n1792_not ; n2999
g2358 and n2998_not n2999_not ; n3000
g2359 and in1[104] n1787 ; n3001
g2360 and in0[104] n1787_not ; n3002
g2361 and n3001_not n3002_not ; n3003
g2362 and n3000_not n3003 ; n3004
g2363 and n2997_not n3004_not ; n3005
g2364 and n2990 n3005 ; n3006
g2365 and n2975_not n3006 ; n3007
g2366 and n2978_not n2981 ; n3008
g2367 and n3000 n3003_not ; n3009
g2368 and n2997_not n3009 ; n3010
g2369 and n2993_not n2996 ; n3011
g2370 and n3010_not n3011_not ; n3012
g2371 and n2985 n2988_not ; n3013
g2372 and n3012 n3013_not ; n3014
g2373 and n2990 n3014_not ; n3015
g2374 and n3008_not n3015_not ; n3016
g2375 and n3007_not n3016 ; n3017
g2376 and n1880 n1883_not ; n3018
g2377 and n1877_not n3018_not ; n3019
g2378 and n1870 n3019 ; n3020
g2379 and n3017_not n3020 ; n3021
g2380 and n1890_not n3021_not ; n3022
g2381 and n1888_not n3022 ; n3023
g2382 and n1861_not n3023 ; n3024
g2383 and n1854_not n3024_not ; n3025
g2384 and n1847 n3025 ; n3026
g2385 and n1832_not n3026 ; n3027
g2386 and n1835_not n1838 ; n3028
g2387 and n1828 n1854_not ; n3029
g2388 and n1831_not n3029 ; n3030
g2389 and n1850_not n1853 ; n3031
g2390 and n3030_not n3031_not ; n3032
g2391 and n1842 n1845_not ; n3033
g2392 and n3032 n3033_not ; n3034
g2393 and n1847 n3034_not ; n3035
g2394 and n3028_not n3035_not ; n3036
g2395 and n3027_not n3036 ; n3037
g2396 and n1808 n1818_not ; n3038
g2397 and n1815_not n3038_not ; n3039
g2398 and n1805 n3039 ; n3040
g2399 and n3037_not n3040 ; n3041
g2400 and n1825_not n3041_not ; n3042
g2401 and n1823_not n3042 ; n3043
g2402 and n1796_not n3043 ; n3044
g2403 and in1[123] n1787 ; n3045
g2404 and in0[123] n1787_not ; n3046
g2405 and n3045_not n3046_not ; n3047
g2406 and in3[123] n1792 ; n3048
g2407 and in2[123] n1792_not ; n3049
g2408 and n3048_not n3049_not ; n3050
g2409 and n3047 n3050_not ; n3051
g2410 and in3[122] n1792 ; n3052
g2411 and in2[122] n1792_not ; n3053
g2412 and n3052_not n3053_not ; n3054
g2413 and in1[122] n1787 ; n3055
g2414 and in0[122] n1787_not ; n3056
g2415 and n3055_not n3056_not ; n3057
g2416 and n3054_not n3057 ; n3058
g2417 and n3051_not n3058_not ; n3059
g2418 and in1[121] n1787 ; n3060
g2419 and in0[121] n1787_not ; n3061
g2420 and n3060_not n3061_not ; n3062
g2421 and in3[121] n1792 ; n3063
g2422 and in2[121] n1792_not ; n3064
g2423 and n3063_not n3064_not ; n3065
g2424 and n3062 n3065_not ; n3066
g2425 and in3[120] n1792 ; n3067
g2426 and in2[120] n1792_not ; n3068
g2427 and n3067_not n3068_not ; n3069
g2428 and in1[120] n1787 ; n3070
g2429 and in0[120] n1787_not ; n3071
g2430 and n3070_not n3071_not ; n3072
g2431 and n3069_not n3072 ; n3073
g2432 and n3066_not n3073_not ; n3074
g2433 and n3059 n3074 ; n3075
g2434 and n3044_not n3075 ; n3076
g2435 and n3047_not n3050 ; n3077
g2436 and n3066_not n3069 ; n3078
g2437 and n3072_not n3078 ; n3079
g2438 and n3062_not n3065 ; n3080
g2439 and n3079_not n3080_not ; n3081
g2440 and n3054 n3057_not ; n3082
g2441 and n3081 n3082_not ; n3083
g2442 and n3059 n3083_not ; n3084
g2443 and n3077_not n3084_not ; n3085
g2444 and n3076_not n3085 ; n3086
g2445 and in1[124] n1787 ; n3087
g2446 and in0[124] n1787_not ; n3088
g2447 and n3087_not n3088_not ; n3089
g2448 and in3[124] n1792 ; n3090
g2449 and in2[124] n1792_not ; n3091
g2450 and n3090_not n3091_not ; n3092
g2451 and n3089 n3092_not ; n3093
g2452 and n1213_not n1784 ; n3094
g2453 and in1[126] n1787 ; n3095
g2454 and in0[126] n1787_not ; n3096
g2455 and n3095_not n3096_not ; n3097
g2456 and in3[126] n1792 ; n3098
g2457 and in2[126] n1792_not ; n3099
g2458 and n3098_not n3099_not ; n3100
g2459 and n3097 n3100_not ; n3101
g2460 and in1[125] n1787 ; n3102
g2461 and in0[125] n1787_not ; n3103
g2462 and n3102_not n3103_not ; n3104
g2463 and in3[125] n1792 ; n3105
g2464 and in2[125] n1792_not ; n3106
g2465 and n3105_not n3106_not ; n3107
g2466 and n3104 n3107_not ; n3108
g2467 and n3101_not n3108_not ; n3109
g2468 and n3094_not n3109 ; n3110
g2469 and n3093_not n3110 ; n3111
g2470 and n3086_not n3111 ; n3112
g2471 and n3089_not n3092 ; n3113
g2472 and n3104_not n3107 ; n3114
g2473 and n3113_not n3114_not ; n3115
g2474 and n3109 n3115_not ; n3116
g2475 and n3097_not n3100 ; n3117
g2476 and n3116_not n3117_not ; n3118
g2477 and n3094_not n3118_not ; n3119
g2478 and n3112_not n3119_not ; n3120
g2479 and n1785_not n3120 ; address[1]
g2480 and n2503_not address[1] ; n3122
g2481 and n2500_not address[1]_not ; n3123
g2482 and n3122_not n3123_not ; result[0]
g2483 and n2497_not address[1] ; n3125
g2484 and n2508_not address[1]_not ; n3126
g2485 and n3125_not n3126_not ; result[1]
g2486 and n2515_not address[1] ; n3128
g2487 and n2512_not address[1]_not ; n3129
g2488 and n3128_not n3129_not ; result[2]
g2489 and n2493_not address[1] ; n3131
g2490 and n2490_not address[1]_not ; n3132
g2491 and n3131_not n3132_not ; result[3]
g2492 and n2484_not address[1] ; n3134
g2493 and n2487_not address[1]_not ; n3135
g2494 and n3134_not n3135_not ; result[4]
g2495 and n2478_not address[1] ; n3137
g2496 and n2481_not address[1]_not ; n3138
g2497 and n3137_not n3138_not ; result[5]
g2498 and n2472_not address[1] ; n3140
g2499 and n2475_not address[1]_not ; n3141
g2500 and n3140_not n3141_not ; result[6]
g2501 and n2468_not address[1] ; n3143
g2502 and n2465_not address[1]_not ; n3144
g2503 and n3143_not n3144_not ; result[7]
g2504 and n2462_not address[1] ; n3146
g2505 and n2542_not address[1]_not ; n3147
g2506 and n3146_not n3147_not ; result[8]
g2507 and n2459_not address[1] ; n3149
g2508 and n2549_not address[1]_not ; n3150
g2509 and n3149_not n3150_not ; result[9]
g2510 and n2455_not address[1] ; n3152
g2511 and n2452_not address[1]_not ; n3153
g2512 and n3152_not n3153_not ; result[10]
g2513 and n2448_not address[1] ; n3155
g2514 and n2445_not address[1]_not ; n3156
g2515 and n3155_not n3156_not ; result[11]
g2516 and n2441_not address[1] ; n3158
g2517 and n2438_not address[1]_not ; n3159
g2518 and n3158_not n3159_not ; result[12]
g2519 and n2434_not address[1] ; n3161
g2520 and n2431_not address[1]_not ; n3162
g2521 and n3161_not n3162_not ; result[13]
g2522 and n2427_not address[1] ; n3164
g2523 and n2424_not address[1]_not ; n3165
g2524 and n3164_not n3165_not ; result[14]
g2525 and n2420_not address[1] ; n3167
g2526 and n2417_not address[1]_not ; n3168
g2527 and n3167_not n3168_not ; result[15]
g2528 and n2414_not address[1] ; n3170
g2529 and n2574_not address[1]_not ; n3171
g2530 and n3170_not n3171_not ; result[16]
g2531 and n2411_not address[1] ; n3173
g2532 and n2581_not address[1]_not ; n3174
g2533 and n3173_not n3174_not ; result[17]
g2534 and n2407_not address[1] ; n3176
g2535 and n2404_not address[1]_not ; n3177
g2536 and n3176_not n3177_not ; result[18]
g2537 and n2400_not address[1] ; n3179
g2538 and n2397_not address[1]_not ; n3180
g2539 and n3179_not n3180_not ; result[19]
g2540 and n2393_not address[1] ; n3182
g2541 and n2390_not address[1]_not ; n3183
g2542 and n3182_not n3183_not ; result[20]
g2543 and n2386_not address[1] ; n3185
g2544 and n2383_not address[1]_not ; n3186
g2545 and n3185_not n3186_not ; result[21]
g2546 and n2379_not address[1] ; n3188
g2547 and n2376_not address[1]_not ; n3189
g2548 and n3188_not n3189_not ; result[22]
g2549 and n2372_not address[1] ; n3191
g2550 and n2369_not address[1]_not ; n3192
g2551 and n3191_not n3192_not ; result[23]
g2552 and n2366_not address[1] ; n3194
g2553 and n2606_not address[1]_not ; n3195
g2554 and n3194_not n3195_not ; result[24]
g2555 and n2363_not address[1] ; n3197
g2556 and n2613_not address[1]_not ; n3198
g2557 and n3197_not n3198_not ; result[25]
g2558 and n2359_not address[1] ; n3200
g2559 and n2356_not address[1]_not ; n3201
g2560 and n3200_not n3201_not ; result[26]
g2561 and n2352_not address[1] ; n3203
g2562 and n2349_not address[1]_not ; n3204
g2563 and n3203_not n3204_not ; result[27]
g2564 and n2345_not address[1] ; n3206
g2565 and n2342_not address[1]_not ; n3207
g2566 and n3206_not n3207_not ; result[28]
g2567 and n2338_not address[1] ; n3209
g2568 and n2335_not address[1]_not ; n3210
g2569 and n3209_not n3210_not ; result[29]
g2570 and n2331_not address[1] ; n3212
g2571 and n2328_not address[1]_not ; n3213
g2572 and n3212_not n3213_not ; result[30]
g2573 and n2324_not address[1] ; n3215
g2574 and n2321_not address[1]_not ; n3216
g2575 and n3215_not n3216_not ; result[31]
g2576 and n2314_not address[1] ; n3218
g2577 and n2317_not address[1]_not ; n3219
g2578 and n3218_not n3219_not ; result[32]
g2579 and n2672_not address[1] ; n3221
g2580 and n2669_not address[1]_not ; n3222
g2581 and n3221_not n3222_not ; result[33]
g2582 and n2683_not address[1] ; n3224
g2583 and n2686_not address[1]_not ; n3225
g2584 and n3224_not n3225_not ; result[34]
g2585 and n2679_not address[1] ; n3227
g2586 and n2676_not address[1]_not ; n3228
g2587 and n3227_not n3228_not ; result[35]
g2588 and n2656_not address[1] ; n3230
g2589 and n2653_not address[1]_not ; n3231
g2590 and n3230_not n3231_not ; result[36]
g2591 and n2663_not address[1] ; n3233
g2592 and n2660_not address[1]_not ; n3234
g2593 and n3233_not n3234_not ; result[37]
g2594 and n2645_not address[1] ; n3236
g2595 and n2648_not address[1]_not ; n3237
g2596 and n3236_not n3237_not ; result[38]
g2597 and n2641_not address[1] ; n3239
g2598 and n2638_not address[1]_not ; n3240
g2599 and n3239_not n3240_not ; result[39]
g2600 and n2295_not address[1] ; n3242
g2601 and n2292_not address[1]_not ; n3243
g2602 and n3242_not n3243_not ; result[40]
g2603 and n2288_not address[1] ; n3245
g2604 and n2285_not address[1]_not ; n3246
g2605 and n3245_not n3246_not ; result[41]
g2606 and n2280_not address[1] ; n3248
g2607 and n2277_not address[1]_not ; n3249
g2608 and n3248_not n3249_not ; result[42]
g2609 and n2272_not address[1] ; n3251
g2610 and n2269_not address[1]_not ; n3252
g2611 and n3251_not n3252_not ; result[43]
g2612 and n2256_not address[1] ; n3254
g2613 and n2253_not address[1]_not ; n3255
g2614 and n3254_not n3255_not ; result[44]
g2615 and n2263_not address[1] ; n3257
g2616 and n2260_not address[1]_not ; n3258
g2617 and n3257_not n3258_not ; result[45]
g2618 and n2245_not address[1] ; n3260
g2619 and n2248_not address[1]_not ; n3261
g2620 and n3260_not n3261_not ; result[46]
g2621 and n2240_not address[1] ; n3263
g2622 and n2237_not address[1]_not ; n3264
g2623 and n3263_not n3264_not ; result[47]
g2624 and n2726_not address[1] ; n3266
g2625 and n2729_not address[1]_not ; n3267
g2626 and n3266_not n3267_not ; result[48]
g2627 and n2767_not address[1] ; n3269
g2628 and n2764_not address[1]_not ; n3270
g2629 and n3269_not n3270_not ; result[49]
g2630 and n2778_not address[1] ; n3272
g2631 and n2781_not address[1]_not ; n3273
g2632 and n3272_not n3273_not ; result[50]
g2633 and n2774_not address[1] ; n3275
g2634 and n2771_not address[1]_not ; n3276
g2635 and n3275_not n3276_not ; result[51]
g2636 and n2755_not address[1] ; n3278
g2637 and n2758_not address[1]_not ; n3279
g2638 and n3278_not n3279_not ; result[52]
g2639 and n2751_not address[1] ; n3281
g2640 and n2748_not address[1]_not ; n3282
g2641 and n3281_not n3282_not ; result[53]
g2642 and n2740_not address[1] ; n3284
g2643 and n2743_not address[1]_not ; n3285
g2644 and n3284_not n3285_not ; result[54]
g2645 and n2736_not address[1] ; n3287
g2646 and n2733_not address[1]_not ; n3288
g2647 and n3287_not n3288_not ; result[55]
g2648 and n2218_not address[1] ; n3290
g2649 and n2215_not address[1]_not ; n3291
g2650 and n3290_not n3291_not ; result[56]
g2651 and n2211_not address[1] ; n3293
g2652 and n2208_not address[1]_not ; n3294
g2653 and n3293_not n3294_not ; result[57]
g2654 and n2203_not address[1] ; n3296
g2655 and n2200_not address[1]_not ; n3297
g2656 and n3296_not n3297_not ; result[58]
g2657 and n2195_not address[1] ; n3299
g2658 and n2192_not address[1]_not ; n3300
g2659 and n3299_not n3300_not ; result[59]
g2660 and n2179_not address[1] ; n3302
g2661 and n2176_not address[1]_not ; n3303
g2662 and n3302_not n3303_not ; result[60]
g2663 and n2186_not address[1] ; n3305
g2664 and n2183_not address[1]_not ; n3306
g2665 and n3305_not n3306_not ; result[61]
g2666 and n2168_not address[1] ; n3308
g2667 and n2171_not address[1]_not ; n3309
g2668 and n3308_not n3309_not ; result[62]
g2669 and n2163_not address[1] ; n3311
g2670 and n2160_not address[1]_not ; n3312
g2671 and n3311_not n3312_not ; result[63]
g2672 and n2146_not address[1] ; n3314
g2673 and n2149_not address[1]_not ; n3315
g2674 and n3314_not n3315_not ; result[64]
g2675 and n2156_not address[1] ; n3317
g2676 and n2153_not address[1]_not ; n3318
g2677 and n3317_not n3318_not ; result[65]
g2678 and n2138_not address[1] ; n3320
g2679 and n2141_not address[1]_not ; n3321
g2680 and n3320_not n3321_not ; result[66]
g2681 and n2134_not address[1] ; n3323
g2682 and n2131_not address[1]_not ; n3324
g2683 and n3323_not n3324_not ; result[67]
g2684 and n2121_not address[1] ; n3326
g2685 and n2118_not address[1]_not ; n3327
g2686 and n3326_not n3327_not ; result[68]
g2687 and n2114_not address[1] ; n3329
g2688 and n2111_not address[1]_not ; n3330
g2689 and n3329_not n3330_not ; result[69]
g2690 and n2103_not address[1] ; n3332
g2691 and n2106_not address[1]_not ; n3333
g2692 and n3332_not n3333_not ; result[70]
g2693 and n2098_not address[1] ; n3335
g2694 and n2095_not address[1]_not ; n3336
g2695 and n3335_not n3336_not ; result[71]
g2696 and n2862_not address[1] ; n3338
g2697 and n2865_not address[1]_not ; n3339
g2698 and n3338_not n3339_not ; result[72]
g2699 and n2858_not address[1] ; n3341
g2700 and n2855_not address[1]_not ; n3342
g2701 and n3341_not n3342_not ; result[73]
g2702 and n2847_not address[1] ; n3344
g2703 and n2850_not address[1]_not ; n3345
g2704 and n3344_not n3345_not ; result[74]
g2705 and n2843_not address[1] ; n3347
g2706 and n2840_not address[1]_not ; n3348
g2707 and n3347_not n3348_not ; result[75]
g2708 and n2085_not address[1] ; n3350
g2709 and n2082_not address[1]_not ; n3351
g2710 and n3350_not n3351_not ; result[76]
g2711 and n2078_not address[1] ; n3353
g2712 and n2075_not address[1]_not ; n3354
g2713 and n3353_not n3354_not ; result[77]
g2714 and n2067_not address[1] ; n3356
g2715 and n2070_not address[1]_not ; n3357
g2716 and n3356_not n3357_not ; result[78]
g2717 and n2062_not address[1] ; n3359
g2718 and n2059_not address[1]_not ; n3360
g2719 and n3359_not n3360_not ; result[79]
g2720 and n2030_not address[1] ; n3362
g2721 and n2033_not address[1]_not ; n3363
g2722 and n3362_not n3363_not ; result[80]
g2723 and n2055_not address[1] ; n3365
g2724 and n2052_not address[1]_not ; n3366
g2725 and n3365_not n3366_not ; result[81]
g2726 and n2044_not address[1] ; n3368
g2727 and n2047_not address[1]_not ; n3369
g2728 and n3368_not n3369_not ; result[82]
g2729 and n2040_not address[1] ; n3371
g2730 and n2037_not address[1]_not ; n3372
g2731 and n3371_not n3372_not ; result[83]
g2732 and n2020_not address[1] ; n3374
g2733 and n2017_not address[1]_not ; n3375
g2734 and n3374_not n3375_not ; result[84]
g2735 and n2013_not address[1] ; n3377
g2736 and n2010_not address[1]_not ; n3378
g2737 and n3377_not n3378_not ; result[85]
g2738 and n2002_not address[1] ; n3380
g2739 and n2005_not address[1]_not ; n3381
g2740 and n3380_not n3381_not ; result[86]
g2741 and n1997_not address[1] ; n3383
g2742 and n1994_not address[1]_not ; n3384
g2743 and n3383_not n3384_not ; result[87]
g2744 and n2931_not address[1] ; n3386
g2745 and n2934_not address[1]_not ; n3387
g2746 and n3386_not n3387_not ; result[88]
g2747 and n2927_not address[1] ; n3389
g2748 and n2924_not address[1]_not ; n3390
g2749 and n3389_not n3390_not ; result[89]
g2750 and n2916_not address[1] ; n3392
g2751 and n2919_not address[1]_not ; n3393
g2752 and n3392_not n3393_not ; result[90]
g2753 and n2912_not address[1] ; n3395
g2754 and n2909_not address[1]_not ; n3396
g2755 and n3395_not n3396_not ; result[91]
g2756 and n1984_not address[1] ; n3398
g2757 and n1981_not address[1]_not ; n3399
g2758 and n3398_not n3399_not ; result[92]
g2759 and n1977_not address[1] ; n3401
g2760 and n1974_not address[1]_not ; n3402
g2761 and n3401_not n3402_not ; result[93]
g2762 and n1966_not address[1] ; n3404
g2763 and n1969_not address[1]_not ; n3405
g2764 and n3404_not n3405_not ; result[94]
g2765 and n1961_not address[1] ; n3407
g2766 and n1958_not address[1]_not ; n3408
g2767 and n3407_not n3408_not ; result[95]
g2768 and n1929_not address[1] ; n3410
g2769 and n1932_not address[1]_not ; n3411
g2770 and n3410_not n3411_not ; result[96]
g2771 and n1954_not address[1] ; n3413
g2772 and n1951_not address[1]_not ; n3414
g2773 and n3413_not n3414_not ; result[97]
g2774 and n1943_not address[1] ; n3416
g2775 and n1946_not address[1]_not ; n3417
g2776 and n3416_not n3417_not ; result[98]
g2777 and n1939_not address[1] ; n3419
g2778 and n1936_not address[1]_not ; n3420
g2779 and n3419_not n3420_not ; result[99]
g2780 and n1919_not address[1] ; n3422
g2781 and n1916_not address[1]_not ; n3423
g2782 and n3422_not n3423_not ; result[100]
g2783 and n1912_not address[1] ; n3425
g2784 and n1909_not address[1]_not ; n3426
g2785 and n3425_not n3426_not ; result[101]
g2786 and n1901_not address[1] ; n3428
g2787 and n1904_not address[1]_not ; n3429
g2788 and n3428_not n3429_not ; result[102]
g2789 and n1896_not address[1] ; n3431
g2790 and n1893_not address[1]_not ; n3432
g2791 and n3431_not n3432_not ; result[103]
g2792 and n3000_not address[1] ; n3434
g2793 and n3003_not address[1]_not ; n3435
g2794 and n3434_not n3435_not ; result[104]
g2795 and n2996_not address[1] ; n3437
g2796 and n2993_not address[1]_not ; n3438
g2797 and n3437_not n3438_not ; result[105]
g2798 and n2985_not address[1] ; n3440
g2799 and n2988_not address[1]_not ; n3441
g2800 and n3440_not n3441_not ; result[106]
g2801 and n2981_not address[1] ; n3443
g2802 and n2978_not address[1]_not ; n3444
g2803 and n3443_not n3444_not ; result[107]
g2804 and n1883_not address[1] ; n3446
g2805 and n1880_not address[1]_not ; n3447
g2806 and n3446_not n3447_not ; result[108]
g2807 and n1876_not address[1] ; n3449
g2808 and n1873_not address[1]_not ; n3450
g2809 and n3449_not n3450_not ; result[109]
g2810 and n1865_not address[1] ; n3452
g2811 and n1868_not address[1]_not ; n3453
g2812 and n3452_not n3453_not ; result[110]
g2813 and n1860_not address[1] ; n3455
g2814 and n1857_not address[1]_not ; n3456
g2815 and n3455_not n3456_not ; result[111]
g2816 and n1828_not address[1] ; n3458
g2817 and n1831_not address[1]_not ; n3459
g2818 and n3458_not n3459_not ; result[112]
g2819 and n1853_not address[1] ; n3461
g2820 and n1850_not address[1]_not ; n3462
g2821 and n3461_not n3462_not ; result[113]
g2822 and n1842_not address[1] ; n3464
g2823 and n1845_not address[1]_not ; n3465
g2824 and n3464_not n3465_not ; result[114]
g2825 and n1838_not address[1] ; n3467
g2826 and n1835_not address[1]_not ; n3468
g2827 and n3467_not n3468_not ; result[115]
g2828 and n1818_not address[1] ; n3470
g2829 and n1808_not address[1]_not ; n3471
g2830 and n3470_not n3471_not ; result[116]
g2831 and n1814_not address[1] ; n3473
g2832 and n1811_not address[1]_not ; n3474
g2833 and n3473_not n3474_not ; result[117]
g2834 and n1800_not address[1] ; n3476
g2835 and n1803_not address[1]_not ; n3477
g2836 and n3476_not n3477_not ; result[118]
g2837 and n1795_not address[1] ; n3479
g2838 and n1790_not address[1]_not ; n3480
g2839 and n3479_not n3480_not ; result[119]
g2840 and n3069_not address[1] ; n3482
g2841 and n3072_not address[1]_not ; n3483
g2842 and n3482_not n3483_not ; result[120]
g2843 and n3065_not address[1] ; n3485
g2844 and n3062_not address[1]_not ; n3486
g2845 and n3485_not n3486_not ; result[121]
g2846 and n3054_not address[1] ; n3488
g2847 and n3057_not address[1]_not ; n3489
g2848 and n3488_not n3489_not ; result[122]
g2849 and n3050_not address[1] ; n3491
g2850 and n3047_not address[1]_not ; n3492
g2851 and n3491_not n3492_not ; result[123]
g2852 and n3092_not address[1] ; n3494
g2853 and n3089_not address[1]_not ; n3495
g2854 and n3494_not n3495_not ; result[124]
g2855 and n3107_not address[1] ; n3497
g2856 and n3104_not address[1]_not ; n3498
g2857 and n3497_not n3498_not ; result[125]
g2858 and n3100_not address[1] ; n3500
g2859 and n3097_not address[1]_not ; n3501
g2860 and n3500_not n3501_not ; result[126]
g2861 and n1213_not n3120 ; n3503
g2862 and n1784 n3503_not ; result[127]
g2863 and n1792 address[1] ; n3505
g2864 and n1787 address[1]_not ; n3506
g2865 and n3505_not n3506_not ; address[0]
g2866 not in3[119] ; in3[119]_not
g2867 not in2[119] ; in2[119]_not
g2868 not in2[118] ; in2[118]_not
g2869 not n644 ; n644_not
g2870 not n645 ; n645_not
g2871 not in2[117] ; in2[117]_not
g2872 not in3[116] ; in3[116]_not
g2873 not n647 ; n647_not
g2874 not in3[117] ; in3[117]_not
g2875 not n649 ; n649_not
g2876 not n650 ; n650_not
g2877 not n651 ; n651_not
g2878 not in3[118] ; in3[118]_not
g2879 not in2[112] ; in2[112]_not
g2880 not in2[115] ; in2[115]_not
g2881 not in2[114] ; in2[114]_not
g2882 not n656 ; n656_not
g2883 not n657 ; n657_not
g2884 not in2[113] ; in2[113]_not
g2885 not in3[111] ; in3[111]_not
g2886 not in2[111] ; in2[111]_not
g2887 not in2[110] ; in2[110]_not
g2888 not n661 ; n661_not
g2889 not n662 ; n662_not
g2890 not in2[109] ; in2[109]_not
g2891 not in3[108] ; in3[108]_not
g2892 not n664 ; n664_not
g2893 not in3[109] ; in3[109]_not
g2894 not n666 ; n666_not
g2895 not n667 ; n667_not
g2896 not n668 ; n668_not
g2897 not in3[110] ; in3[110]_not
g2898 not in3[103] ; in3[103]_not
g2899 not in2[103] ; in2[103]_not
g2900 not in2[102] ; in2[102]_not
g2901 not n673 ; n673_not
g2902 not n674 ; n674_not
g2903 not in2[101] ; in2[101]_not
g2904 not in3[100] ; in3[100]_not
g2905 not n676 ; n676_not
g2906 not in3[101] ; in3[101]_not
g2907 not n678 ; n678_not
g2908 not n679 ; n679_not
g2909 not n680 ; n680_not
g2910 not in3[102] ; in3[102]_not
g2911 not in2[96] ; in2[96]_not
g2912 not in2[99] ; in2[99]_not
g2913 not in2[98] ; in2[98]_not
g2914 not n685 ; n685_not
g2915 not n686 ; n686_not
g2916 not in2[97] ; in2[97]_not
g2917 not in3[95] ; in3[95]_not
g2918 not in2[95] ; in2[95]_not
g2919 not in2[94] ; in2[94]_not
g2920 not n690 ; n690_not
g2921 not n691 ; n691_not
g2922 not in2[93] ; in2[93]_not
g2923 not in3[92] ; in3[92]_not
g2924 not n693 ; n693_not
g2925 not in3[93] ; in3[93]_not
g2926 not n695 ; n695_not
g2927 not n696 ; n696_not
g2928 not n697 ; n697_not
g2929 not in3[94] ; in3[94]_not
g2930 not in3[87] ; in3[87]_not
g2931 not in2[87] ; in2[87]_not
g2932 not in2[86] ; in2[86]_not
g2933 not n702 ; n702_not
g2934 not n703 ; n703_not
g2935 not in2[85] ; in2[85]_not
g2936 not in3[84] ; in3[84]_not
g2937 not n705 ; n705_not
g2938 not in3[85] ; in3[85]_not
g2939 not n707 ; n707_not
g2940 not n708 ; n708_not
g2941 not n709 ; n709_not
g2942 not in3[86] ; in3[86]_not
g2943 not in2[80] ; in2[80]_not
g2944 not in2[83] ; in2[83]_not
g2945 not in2[82] ; in2[82]_not
g2946 not n714 ; n714_not
g2947 not n715 ; n715_not
g2948 not in2[81] ; in2[81]_not
g2949 not in3[79] ; in3[79]_not
g2950 not in2[79] ; in2[79]_not
g2951 not in2[78] ; in2[78]_not
g2952 not n719 ; n719_not
g2953 not n720 ; n720_not
g2954 not in2[77] ; in2[77]_not
g2955 not in3[76] ; in3[76]_not
g2956 not n722 ; n722_not
g2957 not in3[77] ; in3[77]_not
g2958 not n724 ; n724_not
g2959 not n725 ; n725_not
g2960 not n726 ; n726_not
g2961 not in3[78] ; in3[78]_not
g2962 not in3[71] ; in3[71]_not
g2963 not in2[71] ; in2[71]_not
g2964 not in2[70] ; in2[70]_not
g2965 not n731 ; n731_not
g2966 not n732 ; n732_not
g2967 not in2[69] ; in2[69]_not
g2968 not in3[68] ; in3[68]_not
g2969 not n734 ; n734_not
g2970 not in3[69] ; in3[69]_not
g2971 not n736 ; n736_not
g2972 not n737 ; n737_not
g2973 not n738 ; n738_not
g2974 not in3[70] ; in3[70]_not
g2975 not in2[67] ; in2[67]_not
g2976 not in2[66] ; in2[66]_not
g2977 not n742 ; n742_not
g2978 not n743 ; n743_not
g2979 not in2[65] ; in2[65]_not
g2980 not in3[63] ; in3[63]_not
g2981 not in2[63] ; in2[63]_not
g2982 not in2[62] ; in2[62]_not
g2983 not n747 ; n747_not
g2984 not n748 ; n748_not
g2985 not in2[60] ; in2[60]_not
g2986 not in2[61] ; in2[61]_not
g2987 not n750 ; n750_not
g2988 not n751 ; n751_not
g2989 not in3[59] ; in3[59]_not
g2990 not in2[59] ; in2[59]_not
g2991 not in2[58] ; in2[58]_not
g2992 not n755 ; n755_not
g2993 not n756 ; n756_not
g2994 not in2[57] ; in2[57]_not
g2995 not in3[56] ; in3[56]_not
g2996 not n758 ; n758_not
g2997 not in3[57] ; in3[57]_not
g2998 not n760 ; n760_not
g2999 not n761 ; n761_not
g3000 not in3[58] ; in3[58]_not
g3001 not n763 ; n763_not
g3002 not n764 ; n764_not
g3003 not n754 ; n754_not
g3004 not n765 ; n765_not
g3005 not n766 ; n766_not
g3006 not in3[60] ; in3[60]_not
g3007 not in3[61] ; in3[61]_not
g3008 not n769 ; n769_not
g3009 not n770 ; n770_not
g3010 not n771 ; n771_not
g3011 not in3[62] ; in3[62]_not
g3012 not in3[47] ; in3[47]_not
g3013 not in2[47] ; in2[47]_not
g3014 not in2[46] ; in2[46]_not
g3015 not n776 ; n776_not
g3016 not n777 ; n777_not
g3017 not in2[44] ; in2[44]_not
g3018 not in2[45] ; in2[45]_not
g3019 not n779 ; n779_not
g3020 not n780 ; n780_not
g3021 not in3[43] ; in3[43]_not
g3022 not in2[43] ; in2[43]_not
g3023 not in2[42] ; in2[42]_not
g3024 not n784 ; n784_not
g3025 not n785 ; n785_not
g3026 not in2[41] ; in2[41]_not
g3027 not in3[40] ; in3[40]_not
g3028 not n787 ; n787_not
g3029 not in3[41] ; in3[41]_not
g3030 not n789 ; n789_not
g3031 not n790 ; n790_not
g3032 not in3[42] ; in3[42]_not
g3033 not n792 ; n792_not
g3034 not n793 ; n793_not
g3035 not n783 ; n783_not
g3036 not n794 ; n794_not
g3037 not n795 ; n795_not
g3038 not in3[44] ; in3[44]_not
g3039 not in3[45] ; in3[45]_not
g3040 not n798 ; n798_not
g3041 not n799 ; n799_not
g3042 not n800 ; n800_not
g3043 not in3[46] ; in3[46]_not
g3044 not in2[32] ; in2[32]_not
g3045 not in2[31] ; in2[31]_not
g3046 not in2[30] ; in2[30]_not
g3047 not in2[29] ; in2[29]_not
g3048 not in2[28] ; in2[28]_not
g3049 not in2[27] ; in2[27]_not
g3050 not in2[26] ; in2[26]_not
g3051 not in2[23] ; in2[23]_not
g3052 not in2[22] ; in2[22]_not
g3053 not in2[21] ; in2[21]_not
g3054 not in2[20] ; in2[20]_not
g3055 not in2[19] ; in2[19]_not
g3056 not in2[18] ; in2[18]_not
g3057 not in2[15] ; in2[15]_not
g3058 not in2[14] ; in2[14]_not
g3059 not in2[13] ; in2[13]_not
g3060 not in2[12] ; in2[12]_not
g3061 not in2[11] ; in2[11]_not
g3062 not in2[10] ; in2[10]_not
g3063 not in2[7] ; in2[7]_not
g3064 not in2[6] ; in2[6]_not
g3065 not in2[3] ; in2[3]_not
g3066 not in3[0] ; in3[0]_not
g3067 not n827 ; n827_not
g3068 not in2[2] ; in2[2]_not
g3069 not in2[1] ; in2[1]_not
g3070 not n826 ; n826_not
g3071 not n829 ; n829_not
g3072 not n830 ; n830_not
g3073 not n828 ; n828_not
g3074 not in3[2] ; in3[2]_not
g3075 not n832 ; n832_not
g3076 not n833 ; n833_not
g3077 not n825 ; n825_not
g3078 not n834 ; n834_not
g3079 not in3[3] ; in3[3]_not
g3080 not n835 ; n835_not
g3081 not n836 ; n836_not
g3082 not in2[4] ; in2[4]_not
g3083 not in3[4] ; in3[4]_not
g3084 not n838 ; n838_not
g3085 not n837 ; n837_not
g3086 not n839 ; n839_not
g3087 not n840 ; n840_not
g3088 not in2[5] ; in2[5]_not
g3089 not in3[5] ; in3[5]_not
g3090 not n842 ; n842_not
g3091 not n841 ; n841_not
g3092 not n843 ; n843_not
g3093 not n844 ; n844_not
g3094 not n824 ; n824_not
g3095 not n845 ; n845_not
g3096 not in3[6] ; in3[6]_not
g3097 not n846 ; n846_not
g3098 not n847 ; n847_not
g3099 not n823 ; n823_not
g3100 not n848 ; n848_not
g3101 not in3[7] ; in3[7]_not
g3102 not n849 ; n849_not
g3103 not n850 ; n850_not
g3104 not in2[8] ; in2[8]_not
g3105 not in3[8] ; in3[8]_not
g3106 not n852 ; n852_not
g3107 not n851 ; n851_not
g3108 not n853 ; n853_not
g3109 not n854 ; n854_not
g3110 not in2[9] ; in2[9]_not
g3111 not in3[9] ; in3[9]_not
g3112 not n856 ; n856_not
g3113 not n855 ; n855_not
g3114 not n857 ; n857_not
g3115 not n858 ; n858_not
g3116 not n822 ; n822_not
g3117 not n859 ; n859_not
g3118 not in3[10] ; in3[10]_not
g3119 not n860 ; n860_not
g3120 not n861 ; n861_not
g3121 not n821 ; n821_not
g3122 not n862 ; n862_not
g3123 not in3[11] ; in3[11]_not
g3124 not n863 ; n863_not
g3125 not n864 ; n864_not
g3126 not n820 ; n820_not
g3127 not n865 ; n865_not
g3128 not in3[12] ; in3[12]_not
g3129 not n866 ; n866_not
g3130 not n867 ; n867_not
g3131 not n819 ; n819_not
g3132 not n868 ; n868_not
g3133 not in3[13] ; in3[13]_not
g3134 not n869 ; n869_not
g3135 not n870 ; n870_not
g3136 not n818 ; n818_not
g3137 not n871 ; n871_not
g3138 not in3[14] ; in3[14]_not
g3139 not n872 ; n872_not
g3140 not n873 ; n873_not
g3141 not n817 ; n817_not
g3142 not n874 ; n874_not
g3143 not in3[15] ; in3[15]_not
g3144 not n875 ; n875_not
g3145 not n876 ; n876_not
g3146 not in2[16] ; in2[16]_not
g3147 not in3[16] ; in3[16]_not
g3148 not n878 ; n878_not
g3149 not n877 ; n877_not
g3150 not n879 ; n879_not
g3151 not n880 ; n880_not
g3152 not in2[17] ; in2[17]_not
g3153 not in3[17] ; in3[17]_not
g3154 not n882 ; n882_not
g3155 not n881 ; n881_not
g3156 not n883 ; n883_not
g3157 not n884 ; n884_not
g3158 not n816 ; n816_not
g3159 not n885 ; n885_not
g3160 not in3[18] ; in3[18]_not
g3161 not n886 ; n886_not
g3162 not n887 ; n887_not
g3163 not n815 ; n815_not
g3164 not n888 ; n888_not
g3165 not in3[19] ; in3[19]_not
g3166 not n889 ; n889_not
g3167 not n890 ; n890_not
g3168 not n814 ; n814_not
g3169 not n891 ; n891_not
g3170 not in3[20] ; in3[20]_not
g3171 not n892 ; n892_not
g3172 not n893 ; n893_not
g3173 not n813 ; n813_not
g3174 not n894 ; n894_not
g3175 not in3[21] ; in3[21]_not
g3176 not n895 ; n895_not
g3177 not n896 ; n896_not
g3178 not n812 ; n812_not
g3179 not n897 ; n897_not
g3180 not in3[22] ; in3[22]_not
g3181 not n898 ; n898_not
g3182 not n899 ; n899_not
g3183 not n811 ; n811_not
g3184 not n900 ; n900_not
g3185 not in3[23] ; in3[23]_not
g3186 not n901 ; n901_not
g3187 not n902 ; n902_not
g3188 not in2[24] ; in2[24]_not
g3189 not in3[24] ; in3[24]_not
g3190 not n904 ; n904_not
g3191 not n903 ; n903_not
g3192 not n905 ; n905_not
g3193 not n906 ; n906_not
g3194 not in2[25] ; in2[25]_not
g3195 not in3[25] ; in3[25]_not
g3196 not n908 ; n908_not
g3197 not n907 ; n907_not
g3198 not n909 ; n909_not
g3199 not n910 ; n910_not
g3200 not n810 ; n810_not
g3201 not n911 ; n911_not
g3202 not in3[26] ; in3[26]_not
g3203 not n912 ; n912_not
g3204 not n913 ; n913_not
g3205 not n809 ; n809_not
g3206 not n914 ; n914_not
g3207 not in3[27] ; in3[27]_not
g3208 not n915 ; n915_not
g3209 not n916 ; n916_not
g3210 not n808 ; n808_not
g3211 not n917 ; n917_not
g3212 not in3[28] ; in3[28]_not
g3213 not n918 ; n918_not
g3214 not n919 ; n919_not
g3215 not n807 ; n807_not
g3216 not n920 ; n920_not
g3217 not in3[29] ; in3[29]_not
g3218 not n921 ; n921_not
g3219 not n922 ; n922_not
g3220 not n806 ; n806_not
g3221 not n923 ; n923_not
g3222 not in3[30] ; in3[30]_not
g3223 not n924 ; n924_not
g3224 not n925 ; n925_not
g3225 not n805 ; n805_not
g3226 not n926 ; n926_not
g3227 not in3[31] ; in3[31]_not
g3228 not n927 ; n927_not
g3229 not n928 ; n928_not
g3230 not in2[39] ; in2[39]_not
g3231 not in2[38] ; in2[38]_not
g3232 not n930 ; n930_not
g3233 not n931 ; n931_not
g3234 not in2[36] ; in2[36]_not
g3235 not in2[37] ; in2[37]_not
g3236 not n933 ; n933_not
g3237 not n934 ; n934_not
g3238 not in2[33] ; in2[33]_not
g3239 not in2[35] ; in2[35]_not
g3240 not in2[34] ; in2[34]_not
g3241 not n938 ; n938_not
g3242 not n939 ; n939_not
g3243 not n937 ; n937_not
g3244 not n929 ; n929_not
g3245 not n804 ; n804_not
g3246 not in3[39] ; in3[39]_not
g3247 not in3[36] ; in3[36]_not
g3248 not in3[37] ; in3[37]_not
g3249 not n947 ; n947_not
g3250 not n948 ; n948_not
g3251 not n949 ; n949_not
g3252 not in3[38] ; in3[38]_not
g3253 not in3[35] ; in3[35]_not
g3254 not in3[32] ; in3[32]_not
g3255 not in3[33] ; in3[33]_not
g3256 not n955 ; n955_not
g3257 not n956 ; n956_not
g3258 not in3[34] ; in3[34]_not
g3259 not n958 ; n958_not
g3260 not n959 ; n959_not
g3261 not n953 ; n953_not
g3262 not n960 ; n960_not
g3263 not n961 ; n961_not
g3264 not n952 ; n952_not
g3265 not n962 ; n962_not
g3266 not n950 ; n950_not
g3267 not n945 ; n945_not
g3268 not n944 ; n944_not
g3269 not in2[40] ; in2[40]_not
g3270 not n967 ; n967_not
g3271 not n966 ; n966_not
g3272 not n803 ; n803_not
g3273 not n971 ; n971_not
g3274 not n801 ; n801_not
g3275 not n796 ; n796_not
g3276 not n775 ; n775_not
g3277 not in2[48] ; in2[48]_not
g3278 not in2[55] ; in2[55]_not
g3279 not in2[54] ; in2[54]_not
g3280 not n977 ; n977_not
g3281 not n978 ; n978_not
g3282 not in2[53] ; in2[53]_not
g3283 not in2[52] ; in2[52]_not
g3284 not n980 ; n980_not
g3285 not n981 ; n981_not
g3286 not in2[49] ; in2[49]_not
g3287 not in2[51] ; in2[51]_not
g3288 not in2[50] ; in2[50]_not
g3289 not n985 ; n985_not
g3290 not n986 ; n986_not
g3291 not n984 ; n984_not
g3292 not n976 ; n976_not
g3293 not n975 ; n975_not
g3294 not in3[55] ; in3[55]_not
g3295 not in3[51] ; in3[51]_not
g3296 not in3[48] ; in3[48]_not
g3297 not in3[49] ; in3[49]_not
g3298 not n995 ; n995_not
g3299 not n996 ; n996_not
g3300 not in3[50] ; in3[50]_not
g3301 not n998 ; n998_not
g3302 not n999 ; n999_not
g3303 not n993 ; n993_not
g3304 not n1000 ; n1000_not
g3305 not n1001 ; n1001_not
g3306 not in3[52] ; in3[52]_not
g3307 not in3[53] ; in3[53]_not
g3308 not n1004 ; n1004_not
g3309 not n1005 ; n1005_not
g3310 not in3[54] ; in3[54]_not
g3311 not n1007 ; n1007_not
g3312 not n1008 ; n1008_not
g3313 not n1002 ; n1002_not
g3314 not n1009 ; n1009_not
g3315 not n992 ; n992_not
g3316 not n991 ; n991_not
g3317 not in2[56] ; in2[56]_not
g3318 not n1013 ; n1013_not
g3319 not n1012 ; n1012_not
g3320 not n774 ; n774_not
g3321 not n1017 ; n1017_not
g3322 not n772 ; n772_not
g3323 not n767 ; n767_not
g3324 not n746 ; n746_not
g3325 not in2[64] ; in2[64]_not
g3326 not n1021 ; n1021_not
g3327 not n1022 ; n1022_not
g3328 not n745 ; n745_not
g3329 not in3[67] ; in3[67]_not
g3330 not in3[64] ; in3[64]_not
g3331 not in3[65] ; in3[65]_not
g3332 not n1028 ; n1028_not
g3333 not n1029 ; n1029_not
g3334 not in3[66] ; in3[66]_not
g3335 not n1031 ; n1031_not
g3336 not n1032 ; n1032_not
g3337 not n1026 ; n1026_not
g3338 not n1033 ; n1033_not
g3339 not n1025 ; n1025_not
g3340 not in2[68] ; in2[68]_not
g3341 not n1036 ; n1036_not
g3342 not n1035 ; n1035_not
g3343 not n741 ; n741_not
g3344 not n1039 ; n1039_not
g3345 not n739 ; n739_not
g3346 not n730 ; n730_not
g3347 not in2[75] ; in2[75]_not
g3348 not in2[74] ; in2[74]_not
g3349 not n1043 ; n1043_not
g3350 not n1044 ; n1044_not
g3351 not in2[73] ; in2[73]_not
g3352 not in2[72] ; in2[72]_not
g3353 not n1046 ; n1046_not
g3354 not n1047 ; n1047_not
g3355 not n1042 ; n1042_not
g3356 not in3[75] ; in3[75]_not
g3357 not in3[72] ; in3[72]_not
g3358 not in3[73] ; in3[73]_not
g3359 not n1053 ; n1053_not
g3360 not n1054 ; n1054_not
g3361 not in3[74] ; in3[74]_not
g3362 not n1056 ; n1056_not
g3363 not n1057 ; n1057_not
g3364 not n1051 ; n1051_not
g3365 not n1058 ; n1058_not
g3366 not n1050 ; n1050_not
g3367 not in2[76] ; in2[76]_not
g3368 not n1061 ; n1061_not
g3369 not n1060 ; n1060_not
g3370 not n729 ; n729_not
g3371 not n1064 ; n1064_not
g3372 not n727 ; n727_not
g3373 not n718 ; n718_not
g3374 not n717 ; n717_not
g3375 not n1067 ; n1067_not
g3376 not n713 ; n713_not
g3377 not in3[83] ; in3[83]_not
g3378 not in3[80] ; in3[80]_not
g3379 not in3[81] ; in3[81]_not
g3380 not n1073 ; n1073_not
g3381 not n1074 ; n1074_not
g3382 not in3[82] ; in3[82]_not
g3383 not n1076 ; n1076_not
g3384 not n1077 ; n1077_not
g3385 not n1071 ; n1071_not
g3386 not n1078 ; n1078_not
g3387 not n1070 ; n1070_not
g3388 not in2[84] ; in2[84]_not
g3389 not n1081 ; n1081_not
g3390 not n1080 ; n1080_not
g3391 not n712 ; n712_not
g3392 not n1084 ; n1084_not
g3393 not n710 ; n710_not
g3394 not n701 ; n701_not
g3395 not in2[91] ; in2[91]_not
g3396 not in2[90] ; in2[90]_not
g3397 not n1088 ; n1088_not
g3398 not n1089 ; n1089_not
g3399 not in2[89] ; in2[89]_not
g3400 not in2[88] ; in2[88]_not
g3401 not n1091 ; n1091_not
g3402 not n1092 ; n1092_not
g3403 not n1087 ; n1087_not
g3404 not in3[91] ; in3[91]_not
g3405 not in3[88] ; in3[88]_not
g3406 not in3[89] ; in3[89]_not
g3407 not n1098 ; n1098_not
g3408 not n1099 ; n1099_not
g3409 not in3[90] ; in3[90]_not
g3410 not n1101 ; n1101_not
g3411 not n1102 ; n1102_not
g3412 not n1096 ; n1096_not
g3413 not n1103 ; n1103_not
g3414 not n1095 ; n1095_not
g3415 not in2[92] ; in2[92]_not
g3416 not n1106 ; n1106_not
g3417 not n1105 ; n1105_not
g3418 not n700 ; n700_not
g3419 not n1109 ; n1109_not
g3420 not n698 ; n698_not
g3421 not n689 ; n689_not
g3422 not n688 ; n688_not
g3423 not n1112 ; n1112_not
g3424 not n684 ; n684_not
g3425 not in3[99] ; in3[99]_not
g3426 not in3[96] ; in3[96]_not
g3427 not in3[97] ; in3[97]_not
g3428 not n1118 ; n1118_not
g3429 not n1119 ; n1119_not
g3430 not in3[98] ; in3[98]_not
g3431 not n1121 ; n1121_not
g3432 not n1122 ; n1122_not
g3433 not n1116 ; n1116_not
g3434 not n1123 ; n1123_not
g3435 not n1115 ; n1115_not
g3436 not in2[100] ; in2[100]_not
g3437 not n1126 ; n1126_not
g3438 not n1125 ; n1125_not
g3439 not n683 ; n683_not
g3440 not n1129 ; n1129_not
g3441 not n681 ; n681_not
g3442 not n672 ; n672_not
g3443 not in2[107] ; in2[107]_not
g3444 not in2[106] ; in2[106]_not
g3445 not n1133 ; n1133_not
g3446 not n1134 ; n1134_not
g3447 not in2[105] ; in2[105]_not
g3448 not in2[104] ; in2[104]_not
g3449 not n1136 ; n1136_not
g3450 not n1137 ; n1137_not
g3451 not n1132 ; n1132_not
g3452 not in3[107] ; in3[107]_not
g3453 not in3[104] ; in3[104]_not
g3454 not in3[105] ; in3[105]_not
g3455 not n1143 ; n1143_not
g3456 not n1144 ; n1144_not
g3457 not in3[106] ; in3[106]_not
g3458 not n1146 ; n1146_not
g3459 not n1147 ; n1147_not
g3460 not n1141 ; n1141_not
g3461 not n1148 ; n1148_not
g3462 not n1140 ; n1140_not
g3463 not in2[108] ; in2[108]_not
g3464 not n1151 ; n1151_not
g3465 not n1150 ; n1150_not
g3466 not n671 ; n671_not
g3467 not n1154 ; n1154_not
g3468 not n669 ; n669_not
g3469 not n660 ; n660_not
g3470 not n659 ; n659_not
g3471 not n1157 ; n1157_not
g3472 not n655 ; n655_not
g3473 not in3[115] ; in3[115]_not
g3474 not in3[112] ; in3[112]_not
g3475 not in3[113] ; in3[113]_not
g3476 not n1163 ; n1163_not
g3477 not n1164 ; n1164_not
g3478 not in3[114] ; in3[114]_not
g3479 not n1166 ; n1166_not
g3480 not n1167 ; n1167_not
g3481 not n1161 ; n1161_not
g3482 not n1168 ; n1168_not
g3483 not n1160 ; n1160_not
g3484 not in2[116] ; in2[116]_not
g3485 not n1171 ; n1171_not
g3486 not n1170 ; n1170_not
g3487 not n654 ; n654_not
g3488 not n1174 ; n1174_not
g3489 not n652 ; n652_not
g3490 not n643 ; n643_not
g3491 not in2[123] ; in2[123]_not
g3492 not in2[122] ; in2[122]_not
g3493 not n1178 ; n1178_not
g3494 not n1179 ; n1179_not
g3495 not in2[121] ; in2[121]_not
g3496 not in2[120] ; in2[120]_not
g3497 not n1181 ; n1181_not
g3498 not n1182 ; n1182_not
g3499 not n1177 ; n1177_not
g3500 not in3[123] ; in3[123]_not
g3501 not in3[120] ; in3[120]_not
g3502 not in3[121] ; in3[121]_not
g3503 not n1188 ; n1188_not
g3504 not n1189 ; n1189_not
g3505 not in3[122] ; in3[122]_not
g3506 not n1191 ; n1191_not
g3507 not n1192 ; n1192_not
g3508 not n1186 ; n1186_not
g3509 not n1193 ; n1193_not
g3510 not n1185 ; n1185_not
g3511 not in2[124] ; in2[124]_not
g3512 not in3[127] ; in3[127]_not
g3513 not in2[126] ; in2[126]_not
g3514 not in2[125] ; in2[125]_not
g3515 not n1198 ; n1198_not
g3516 not n1199 ; n1199_not
g3517 not n1197 ; n1197_not
g3518 not n1196 ; n1196_not
g3519 not n1195 ; n1195_not
g3520 not in3[124] ; in3[124]_not
g3521 not in3[125] ; in3[125]_not
g3522 not n1204 ; n1204_not
g3523 not n1205 ; n1205_not
g3524 not n1206 ; n1206_not
g3525 not in3[126] ; in3[126]_not
g3526 not n1207 ; n1207_not
g3527 not n1208 ; n1208_not
g3528 not n1209 ; n1209_not
g3529 not n1203 ; n1203_not
g3530 not n1210 ; n1210_not
g3531 not n1212 ; n1212_not
g3532 not in1[119] ; in1[119]_not
g3533 not in0[119] ; in0[119]_not
g3534 not in0[118] ; in0[118]_not
g3535 not n1215 ; n1215_not
g3536 not n1216 ; n1216_not
g3537 not in0[117] ; in0[117]_not
g3538 not in1[116] ; in1[116]_not
g3539 not n1218 ; n1218_not
g3540 not in1[117] ; in1[117]_not
g3541 not n1220 ; n1220_not
g3542 not n1221 ; n1221_not
g3543 not n1222 ; n1222_not
g3544 not in1[118] ; in1[118]_not
g3545 not in0[112] ; in0[112]_not
g3546 not in0[115] ; in0[115]_not
g3547 not in0[114] ; in0[114]_not
g3548 not n1227 ; n1227_not
g3549 not n1228 ; n1228_not
g3550 not in0[113] ; in0[113]_not
g3551 not in1[111] ; in1[111]_not
g3552 not in0[111] ; in0[111]_not
g3553 not in0[110] ; in0[110]_not
g3554 not n1232 ; n1232_not
g3555 not n1233 ; n1233_not
g3556 not in0[109] ; in0[109]_not
g3557 not in1[108] ; in1[108]_not
g3558 not n1235 ; n1235_not
g3559 not in1[109] ; in1[109]_not
g3560 not n1237 ; n1237_not
g3561 not n1238 ; n1238_not
g3562 not n1239 ; n1239_not
g3563 not in1[110] ; in1[110]_not
g3564 not in1[103] ; in1[103]_not
g3565 not in0[103] ; in0[103]_not
g3566 not in0[102] ; in0[102]_not
g3567 not n1244 ; n1244_not
g3568 not n1245 ; n1245_not
g3569 not in0[101] ; in0[101]_not
g3570 not in1[100] ; in1[100]_not
g3571 not n1247 ; n1247_not
g3572 not in1[101] ; in1[101]_not
g3573 not n1249 ; n1249_not
g3574 not n1250 ; n1250_not
g3575 not n1251 ; n1251_not
g3576 not in1[102] ; in1[102]_not
g3577 not in0[96] ; in0[96]_not
g3578 not in0[99] ; in0[99]_not
g3579 not in0[98] ; in0[98]_not
g3580 not n1256 ; n1256_not
g3581 not n1257 ; n1257_not
g3582 not in0[97] ; in0[97]_not
g3583 not in1[95] ; in1[95]_not
g3584 not in0[95] ; in0[95]_not
g3585 not in0[94] ; in0[94]_not
g3586 not n1261 ; n1261_not
g3587 not n1262 ; n1262_not
g3588 not in0[93] ; in0[93]_not
g3589 not in1[92] ; in1[92]_not
g3590 not n1264 ; n1264_not
g3591 not in1[93] ; in1[93]_not
g3592 not n1266 ; n1266_not
g3593 not n1267 ; n1267_not
g3594 not n1268 ; n1268_not
g3595 not in1[94] ; in1[94]_not
g3596 not in1[87] ; in1[87]_not
g3597 not in0[87] ; in0[87]_not
g3598 not in0[86] ; in0[86]_not
g3599 not n1273 ; n1273_not
g3600 not n1274 ; n1274_not
g3601 not in0[85] ; in0[85]_not
g3602 not in1[84] ; in1[84]_not
g3603 not n1276 ; n1276_not
g3604 not in1[85] ; in1[85]_not
g3605 not n1278 ; n1278_not
g3606 not n1279 ; n1279_not
g3607 not n1280 ; n1280_not
g3608 not in1[86] ; in1[86]_not
g3609 not in0[80] ; in0[80]_not
g3610 not in0[83] ; in0[83]_not
g3611 not in0[82] ; in0[82]_not
g3612 not n1285 ; n1285_not
g3613 not n1286 ; n1286_not
g3614 not in0[81] ; in0[81]_not
g3615 not in1[79] ; in1[79]_not
g3616 not in0[79] ; in0[79]_not
g3617 not in0[78] ; in0[78]_not
g3618 not n1290 ; n1290_not
g3619 not n1291 ; n1291_not
g3620 not in0[77] ; in0[77]_not
g3621 not in1[76] ; in1[76]_not
g3622 not n1293 ; n1293_not
g3623 not in1[77] ; in1[77]_not
g3624 not n1295 ; n1295_not
g3625 not n1296 ; n1296_not
g3626 not n1297 ; n1297_not
g3627 not in1[78] ; in1[78]_not
g3628 not in1[71] ; in1[71]_not
g3629 not in0[71] ; in0[71]_not
g3630 not in0[70] ; in0[70]_not
g3631 not n1302 ; n1302_not
g3632 not n1303 ; n1303_not
g3633 not in0[69] ; in0[69]_not
g3634 not in1[68] ; in1[68]_not
g3635 not n1305 ; n1305_not
g3636 not in1[69] ; in1[69]_not
g3637 not n1307 ; n1307_not
g3638 not n1308 ; n1308_not
g3639 not n1309 ; n1309_not
g3640 not in1[70] ; in1[70]_not
g3641 not in0[67] ; in0[67]_not
g3642 not in0[66] ; in0[66]_not
g3643 not n1313 ; n1313_not
g3644 not n1314 ; n1314_not
g3645 not in0[65] ; in0[65]_not
g3646 not in1[63] ; in1[63]_not
g3647 not in0[63] ; in0[63]_not
g3648 not in0[62] ; in0[62]_not
g3649 not n1318 ; n1318_not
g3650 not n1319 ; n1319_not
g3651 not in0[60] ; in0[60]_not
g3652 not in0[61] ; in0[61]_not
g3653 not n1321 ; n1321_not
g3654 not n1322 ; n1322_not
g3655 not in1[59] ; in1[59]_not
g3656 not in0[59] ; in0[59]_not
g3657 not in0[58] ; in0[58]_not
g3658 not n1326 ; n1326_not
g3659 not n1327 ; n1327_not
g3660 not in0[57] ; in0[57]_not
g3661 not in1[56] ; in1[56]_not
g3662 not n1329 ; n1329_not
g3663 not in1[57] ; in1[57]_not
g3664 not n1331 ; n1331_not
g3665 not n1332 ; n1332_not
g3666 not in1[58] ; in1[58]_not
g3667 not n1334 ; n1334_not
g3668 not n1335 ; n1335_not
g3669 not n1325 ; n1325_not
g3670 not n1336 ; n1336_not
g3671 not n1337 ; n1337_not
g3672 not in1[60] ; in1[60]_not
g3673 not in1[61] ; in1[61]_not
g3674 not n1340 ; n1340_not
g3675 not n1341 ; n1341_not
g3676 not n1342 ; n1342_not
g3677 not in1[62] ; in1[62]_not
g3678 not in1[47] ; in1[47]_not
g3679 not in0[47] ; in0[47]_not
g3680 not in0[46] ; in0[46]_not
g3681 not n1347 ; n1347_not
g3682 not n1348 ; n1348_not
g3683 not in0[44] ; in0[44]_not
g3684 not in0[45] ; in0[45]_not
g3685 not n1350 ; n1350_not
g3686 not n1351 ; n1351_not
g3687 not in1[43] ; in1[43]_not
g3688 not in0[43] ; in0[43]_not
g3689 not in0[42] ; in0[42]_not
g3690 not n1355 ; n1355_not
g3691 not n1356 ; n1356_not
g3692 not in0[41] ; in0[41]_not
g3693 not in1[40] ; in1[40]_not
g3694 not n1358 ; n1358_not
g3695 not in1[41] ; in1[41]_not
g3696 not n1360 ; n1360_not
g3697 not n1361 ; n1361_not
g3698 not in1[42] ; in1[42]_not
g3699 not n1363 ; n1363_not
g3700 not n1364 ; n1364_not
g3701 not n1354 ; n1354_not
g3702 not n1365 ; n1365_not
g3703 not n1366 ; n1366_not
g3704 not in1[44] ; in1[44]_not
g3705 not in1[45] ; in1[45]_not
g3706 not n1369 ; n1369_not
g3707 not n1370 ; n1370_not
g3708 not n1371 ; n1371_not
g3709 not in1[46] ; in1[46]_not
g3710 not in0[32] ; in0[32]_not
g3711 not in0[31] ; in0[31]_not
g3712 not in0[30] ; in0[30]_not
g3713 not in0[29] ; in0[29]_not
g3714 not in0[28] ; in0[28]_not
g3715 not in0[27] ; in0[27]_not
g3716 not in0[26] ; in0[26]_not
g3717 not in0[23] ; in0[23]_not
g3718 not in0[22] ; in0[22]_not
g3719 not in0[21] ; in0[21]_not
g3720 not in0[20] ; in0[20]_not
g3721 not in0[19] ; in0[19]_not
g3722 not in0[18] ; in0[18]_not
g3723 not in0[15] ; in0[15]_not
g3724 not in0[14] ; in0[14]_not
g3725 not in0[13] ; in0[13]_not
g3726 not in0[12] ; in0[12]_not
g3727 not in0[11] ; in0[11]_not
g3728 not in0[10] ; in0[10]_not
g3729 not in0[7] ; in0[7]_not
g3730 not in0[6] ; in0[6]_not
g3731 not in0[3] ; in0[3]_not
g3732 not in1[0] ; in1[0]_not
g3733 not in1[1] ; in1[1]_not
g3734 not n1397 ; n1397_not
g3735 not n1398 ; n1398_not
g3736 not in0[2] ; in0[2]_not
g3737 not in0[1] ; in0[1]_not
g3738 not n1400 ; n1400_not
g3739 not n1401 ; n1401_not
g3740 not n1399 ; n1399_not
g3741 not in1[2] ; in1[2]_not
g3742 not n1403 ; n1403_not
g3743 not n1404 ; n1404_not
g3744 not n1396 ; n1396_not
g3745 not n1405 ; n1405_not
g3746 not in1[3] ; in1[3]_not
g3747 not n1406 ; n1406_not
g3748 not n1407 ; n1407_not
g3749 not in0[4] ; in0[4]_not
g3750 not in1[4] ; in1[4]_not
g3751 not n1409 ; n1409_not
g3752 not n1408 ; n1408_not
g3753 not n1410 ; n1410_not
g3754 not n1411 ; n1411_not
g3755 not in0[5] ; in0[5]_not
g3756 not in1[5] ; in1[5]_not
g3757 not n1413 ; n1413_not
g3758 not n1412 ; n1412_not
g3759 not n1414 ; n1414_not
g3760 not n1415 ; n1415_not
g3761 not n1395 ; n1395_not
g3762 not n1416 ; n1416_not
g3763 not in1[6] ; in1[6]_not
g3764 not n1417 ; n1417_not
g3765 not n1418 ; n1418_not
g3766 not n1394 ; n1394_not
g3767 not n1419 ; n1419_not
g3768 not in1[7] ; in1[7]_not
g3769 not n1420 ; n1420_not
g3770 not n1421 ; n1421_not
g3771 not in0[8] ; in0[8]_not
g3772 not in1[8] ; in1[8]_not
g3773 not n1423 ; n1423_not
g3774 not n1422 ; n1422_not
g3775 not n1424 ; n1424_not
g3776 not n1425 ; n1425_not
g3777 not in0[9] ; in0[9]_not
g3778 not in1[9] ; in1[9]_not
g3779 not n1427 ; n1427_not
g3780 not n1426 ; n1426_not
g3781 not n1428 ; n1428_not
g3782 not n1429 ; n1429_not
g3783 not n1393 ; n1393_not
g3784 not n1430 ; n1430_not
g3785 not in1[10] ; in1[10]_not
g3786 not n1431 ; n1431_not
g3787 not n1432 ; n1432_not
g3788 not n1392 ; n1392_not
g3789 not n1433 ; n1433_not
g3790 not in1[11] ; in1[11]_not
g3791 not n1434 ; n1434_not
g3792 not n1435 ; n1435_not
g3793 not n1391 ; n1391_not
g3794 not n1436 ; n1436_not
g3795 not in1[12] ; in1[12]_not
g3796 not n1437 ; n1437_not
g3797 not n1438 ; n1438_not
g3798 not n1390 ; n1390_not
g3799 not n1439 ; n1439_not
g3800 not in1[13] ; in1[13]_not
g3801 not n1440 ; n1440_not
g3802 not n1441 ; n1441_not
g3803 not n1389 ; n1389_not
g3804 not n1442 ; n1442_not
g3805 not in1[14] ; in1[14]_not
g3806 not n1443 ; n1443_not
g3807 not n1444 ; n1444_not
g3808 not n1388 ; n1388_not
g3809 not n1445 ; n1445_not
g3810 not in1[15] ; in1[15]_not
g3811 not n1446 ; n1446_not
g3812 not n1447 ; n1447_not
g3813 not in0[16] ; in0[16]_not
g3814 not in1[16] ; in1[16]_not
g3815 not n1449 ; n1449_not
g3816 not n1448 ; n1448_not
g3817 not n1450 ; n1450_not
g3818 not n1451 ; n1451_not
g3819 not in0[17] ; in0[17]_not
g3820 not in1[17] ; in1[17]_not
g3821 not n1453 ; n1453_not
g3822 not n1452 ; n1452_not
g3823 not n1454 ; n1454_not
g3824 not n1455 ; n1455_not
g3825 not n1387 ; n1387_not
g3826 not n1456 ; n1456_not
g3827 not in1[18] ; in1[18]_not
g3828 not n1457 ; n1457_not
g3829 not n1458 ; n1458_not
g3830 not n1386 ; n1386_not
g3831 not n1459 ; n1459_not
g3832 not in1[19] ; in1[19]_not
g3833 not n1460 ; n1460_not
g3834 not n1461 ; n1461_not
g3835 not n1385 ; n1385_not
g3836 not n1462 ; n1462_not
g3837 not in1[20] ; in1[20]_not
g3838 not n1463 ; n1463_not
g3839 not n1464 ; n1464_not
g3840 not n1384 ; n1384_not
g3841 not n1465 ; n1465_not
g3842 not in1[21] ; in1[21]_not
g3843 not n1466 ; n1466_not
g3844 not n1467 ; n1467_not
g3845 not n1383 ; n1383_not
g3846 not n1468 ; n1468_not
g3847 not in1[22] ; in1[22]_not
g3848 not n1469 ; n1469_not
g3849 not n1470 ; n1470_not
g3850 not n1382 ; n1382_not
g3851 not n1471 ; n1471_not
g3852 not in1[23] ; in1[23]_not
g3853 not n1472 ; n1472_not
g3854 not n1473 ; n1473_not
g3855 not in0[24] ; in0[24]_not
g3856 not in1[24] ; in1[24]_not
g3857 not n1475 ; n1475_not
g3858 not n1474 ; n1474_not
g3859 not n1476 ; n1476_not
g3860 not n1477 ; n1477_not
g3861 not in0[25] ; in0[25]_not
g3862 not in1[25] ; in1[25]_not
g3863 not n1479 ; n1479_not
g3864 not n1478 ; n1478_not
g3865 not n1480 ; n1480_not
g3866 not n1481 ; n1481_not
g3867 not n1381 ; n1381_not
g3868 not n1482 ; n1482_not
g3869 not in1[26] ; in1[26]_not
g3870 not n1483 ; n1483_not
g3871 not n1484 ; n1484_not
g3872 not n1380 ; n1380_not
g3873 not n1485 ; n1485_not
g3874 not in1[27] ; in1[27]_not
g3875 not n1486 ; n1486_not
g3876 not n1487 ; n1487_not
g3877 not n1379 ; n1379_not
g3878 not n1488 ; n1488_not
g3879 not in1[28] ; in1[28]_not
g3880 not n1489 ; n1489_not
g3881 not n1490 ; n1490_not
g3882 not n1378 ; n1378_not
g3883 not n1491 ; n1491_not
g3884 not in1[29] ; in1[29]_not
g3885 not n1492 ; n1492_not
g3886 not n1493 ; n1493_not
g3887 not n1377 ; n1377_not
g3888 not n1494 ; n1494_not
g3889 not in1[30] ; in1[30]_not
g3890 not n1495 ; n1495_not
g3891 not n1496 ; n1496_not
g3892 not n1376 ; n1376_not
g3893 not n1497 ; n1497_not
g3894 not in1[31] ; in1[31]_not
g3895 not n1498 ; n1498_not
g3896 not n1499 ; n1499_not
g3897 not in0[39] ; in0[39]_not
g3898 not in0[38] ; in0[38]_not
g3899 not n1501 ; n1501_not
g3900 not n1502 ; n1502_not
g3901 not in0[36] ; in0[36]_not
g3902 not in0[37] ; in0[37]_not
g3903 not n1504 ; n1504_not
g3904 not n1505 ; n1505_not
g3905 not in0[33] ; in0[33]_not
g3906 not in0[35] ; in0[35]_not
g3907 not in0[34] ; in0[34]_not
g3908 not n1509 ; n1509_not
g3909 not n1510 ; n1510_not
g3910 not n1508 ; n1508_not
g3911 not n1500 ; n1500_not
g3912 not n1375 ; n1375_not
g3913 not in1[39] ; in1[39]_not
g3914 not in1[36] ; in1[36]_not
g3915 not in1[37] ; in1[37]_not
g3916 not n1518 ; n1518_not
g3917 not n1519 ; n1519_not
g3918 not n1520 ; n1520_not
g3919 not in1[38] ; in1[38]_not
g3920 not in1[35] ; in1[35]_not
g3921 not in1[32] ; in1[32]_not
g3922 not in1[33] ; in1[33]_not
g3923 not n1526 ; n1526_not
g3924 not n1527 ; n1527_not
g3925 not in1[34] ; in1[34]_not
g3926 not n1529 ; n1529_not
g3927 not n1530 ; n1530_not
g3928 not n1524 ; n1524_not
g3929 not n1531 ; n1531_not
g3930 not n1532 ; n1532_not
g3931 not n1523 ; n1523_not
g3932 not n1533 ; n1533_not
g3933 not n1521 ; n1521_not
g3934 not n1516 ; n1516_not
g3935 not n1515 ; n1515_not
g3936 not in0[40] ; in0[40]_not
g3937 not n1538 ; n1538_not
g3938 not n1537 ; n1537_not
g3939 not n1374 ; n1374_not
g3940 not n1542 ; n1542_not
g3941 not n1372 ; n1372_not
g3942 not n1367 ; n1367_not
g3943 not n1346 ; n1346_not
g3944 not in0[48] ; in0[48]_not
g3945 not in0[55] ; in0[55]_not
g3946 not in0[54] ; in0[54]_not
g3947 not n1548 ; n1548_not
g3948 not n1549 ; n1549_not
g3949 not in0[53] ; in0[53]_not
g3950 not in0[52] ; in0[52]_not
g3951 not n1551 ; n1551_not
g3952 not n1552 ; n1552_not
g3953 not in0[49] ; in0[49]_not
g3954 not in0[51] ; in0[51]_not
g3955 not in0[50] ; in0[50]_not
g3956 not n1556 ; n1556_not
g3957 not n1557 ; n1557_not
g3958 not n1555 ; n1555_not
g3959 not n1547 ; n1547_not
g3960 not n1546 ; n1546_not
g3961 not in1[55] ; in1[55]_not
g3962 not in1[51] ; in1[51]_not
g3963 not in1[48] ; in1[48]_not
g3964 not in1[49] ; in1[49]_not
g3965 not n1566 ; n1566_not
g3966 not n1567 ; n1567_not
g3967 not in1[50] ; in1[50]_not
g3968 not n1569 ; n1569_not
g3969 not n1570 ; n1570_not
g3970 not n1564 ; n1564_not
g3971 not n1571 ; n1571_not
g3972 not n1572 ; n1572_not
g3973 not in1[52] ; in1[52]_not
g3974 not in1[53] ; in1[53]_not
g3975 not n1575 ; n1575_not
g3976 not n1576 ; n1576_not
g3977 not in1[54] ; in1[54]_not
g3978 not n1578 ; n1578_not
g3979 not n1579 ; n1579_not
g3980 not n1573 ; n1573_not
g3981 not n1580 ; n1580_not
g3982 not n1563 ; n1563_not
g3983 not n1562 ; n1562_not
g3984 not in0[56] ; in0[56]_not
g3985 not n1584 ; n1584_not
g3986 not n1583 ; n1583_not
g3987 not n1345 ; n1345_not
g3988 not n1588 ; n1588_not
g3989 not n1343 ; n1343_not
g3990 not n1338 ; n1338_not
g3991 not n1317 ; n1317_not
g3992 not in0[64] ; in0[64]_not
g3993 not n1592 ; n1592_not
g3994 not n1593 ; n1593_not
g3995 not n1316 ; n1316_not
g3996 not in1[67] ; in1[67]_not
g3997 not in1[64] ; in1[64]_not
g3998 not in1[65] ; in1[65]_not
g3999 not n1599 ; n1599_not
g4000 not n1600 ; n1600_not
g4001 not in1[66] ; in1[66]_not
g4002 not n1602 ; n1602_not
g4003 not n1603 ; n1603_not
g4004 not n1597 ; n1597_not
g4005 not n1604 ; n1604_not
g4006 not n1596 ; n1596_not
g4007 not in0[68] ; in0[68]_not
g4008 not n1607 ; n1607_not
g4009 not n1606 ; n1606_not
g4010 not n1312 ; n1312_not
g4011 not n1610 ; n1610_not
g4012 not n1310 ; n1310_not
g4013 not n1301 ; n1301_not
g4014 not in0[75] ; in0[75]_not
g4015 not in0[74] ; in0[74]_not
g4016 not n1614 ; n1614_not
g4017 not n1615 ; n1615_not
g4018 not in0[73] ; in0[73]_not
g4019 not in0[72] ; in0[72]_not
g4020 not n1617 ; n1617_not
g4021 not n1618 ; n1618_not
g4022 not n1613 ; n1613_not
g4023 not in1[75] ; in1[75]_not
g4024 not in1[72] ; in1[72]_not
g4025 not in1[73] ; in1[73]_not
g4026 not n1624 ; n1624_not
g4027 not n1625 ; n1625_not
g4028 not in1[74] ; in1[74]_not
g4029 not n1627 ; n1627_not
g4030 not n1628 ; n1628_not
g4031 not n1622 ; n1622_not
g4032 not n1629 ; n1629_not
g4033 not n1621 ; n1621_not
g4034 not in0[76] ; in0[76]_not
g4035 not n1632 ; n1632_not
g4036 not n1631 ; n1631_not
g4037 not n1300 ; n1300_not
g4038 not n1635 ; n1635_not
g4039 not n1298 ; n1298_not
g4040 not n1289 ; n1289_not
g4041 not n1288 ; n1288_not
g4042 not n1638 ; n1638_not
g4043 not n1284 ; n1284_not
g4044 not in1[83] ; in1[83]_not
g4045 not in1[80] ; in1[80]_not
g4046 not in1[81] ; in1[81]_not
g4047 not n1644 ; n1644_not
g4048 not n1645 ; n1645_not
g4049 not in1[82] ; in1[82]_not
g4050 not n1647 ; n1647_not
g4051 not n1648 ; n1648_not
g4052 not n1642 ; n1642_not
g4053 not n1649 ; n1649_not
g4054 not n1641 ; n1641_not
g4055 not in0[84] ; in0[84]_not
g4056 not n1652 ; n1652_not
g4057 not n1651 ; n1651_not
g4058 not n1283 ; n1283_not
g4059 not n1655 ; n1655_not
g4060 not n1281 ; n1281_not
g4061 not n1272 ; n1272_not
g4062 not in0[91] ; in0[91]_not
g4063 not in0[90] ; in0[90]_not
g4064 not n1659 ; n1659_not
g4065 not n1660 ; n1660_not
g4066 not in0[89] ; in0[89]_not
g4067 not in0[88] ; in0[88]_not
g4068 not n1662 ; n1662_not
g4069 not n1663 ; n1663_not
g4070 not n1658 ; n1658_not
g4071 not in1[91] ; in1[91]_not
g4072 not in1[88] ; in1[88]_not
g4073 not in1[89] ; in1[89]_not
g4074 not n1669 ; n1669_not
g4075 not n1670 ; n1670_not
g4076 not in1[90] ; in1[90]_not
g4077 not n1672 ; n1672_not
g4078 not n1673 ; n1673_not
g4079 not n1667 ; n1667_not
g4080 not n1674 ; n1674_not
g4081 not n1666 ; n1666_not
g4082 not in0[92] ; in0[92]_not
g4083 not n1677 ; n1677_not
g4084 not n1676 ; n1676_not
g4085 not n1271 ; n1271_not
g4086 not n1680 ; n1680_not
g4087 not n1269 ; n1269_not
g4088 not n1260 ; n1260_not
g4089 not n1259 ; n1259_not
g4090 not n1683 ; n1683_not
g4091 not n1255 ; n1255_not
g4092 not in1[99] ; in1[99]_not
g4093 not in1[96] ; in1[96]_not
g4094 not in1[97] ; in1[97]_not
g4095 not n1689 ; n1689_not
g4096 not n1690 ; n1690_not
g4097 not in1[98] ; in1[98]_not
g4098 not n1692 ; n1692_not
g4099 not n1693 ; n1693_not
g4100 not n1687 ; n1687_not
g4101 not n1694 ; n1694_not
g4102 not n1686 ; n1686_not
g4103 not in0[100] ; in0[100]_not
g4104 not n1697 ; n1697_not
g4105 not n1696 ; n1696_not
g4106 not n1254 ; n1254_not
g4107 not n1700 ; n1700_not
g4108 not n1252 ; n1252_not
g4109 not n1243 ; n1243_not
g4110 not in0[107] ; in0[107]_not
g4111 not in0[106] ; in0[106]_not
g4112 not n1704 ; n1704_not
g4113 not n1705 ; n1705_not
g4114 not in0[105] ; in0[105]_not
g4115 not in0[104] ; in0[104]_not
g4116 not n1707 ; n1707_not
g4117 not n1708 ; n1708_not
g4118 not n1703 ; n1703_not
g4119 not in1[107] ; in1[107]_not
g4120 not in1[104] ; in1[104]_not
g4121 not in1[105] ; in1[105]_not
g4122 not n1714 ; n1714_not
g4123 not n1715 ; n1715_not
g4124 not in1[106] ; in1[106]_not
g4125 not n1717 ; n1717_not
g4126 not n1718 ; n1718_not
g4127 not n1712 ; n1712_not
g4128 not n1719 ; n1719_not
g4129 not n1711 ; n1711_not
g4130 not in0[108] ; in0[108]_not
g4131 not n1722 ; n1722_not
g4132 not n1721 ; n1721_not
g4133 not n1242 ; n1242_not
g4134 not n1725 ; n1725_not
g4135 not n1240 ; n1240_not
g4136 not n1231 ; n1231_not
g4137 not n1230 ; n1230_not
g4138 not n1728 ; n1728_not
g4139 not n1226 ; n1226_not
g4140 not in1[115] ; in1[115]_not
g4141 not in1[112] ; in1[112]_not
g4142 not in1[113] ; in1[113]_not
g4143 not n1734 ; n1734_not
g4144 not n1735 ; n1735_not
g4145 not in1[114] ; in1[114]_not
g4146 not n1737 ; n1737_not
g4147 not n1738 ; n1738_not
g4148 not n1732 ; n1732_not
g4149 not n1739 ; n1739_not
g4150 not n1731 ; n1731_not
g4151 not in0[116] ; in0[116]_not
g4152 not n1742 ; n1742_not
g4153 not n1741 ; n1741_not
g4154 not n1225 ; n1225_not
g4155 not n1745 ; n1745_not
g4156 not n1223 ; n1223_not
g4157 not n1214 ; n1214_not
g4158 not in0[123] ; in0[123]_not
g4159 not in0[122] ; in0[122]_not
g4160 not n1749 ; n1749_not
g4161 not n1750 ; n1750_not
g4162 not in0[121] ; in0[121]_not
g4163 not in0[120] ; in0[120]_not
g4164 not n1752 ; n1752_not
g4165 not n1753 ; n1753_not
g4166 not n1748 ; n1748_not
g4167 not in1[123] ; in1[123]_not
g4168 not in1[120] ; in1[120]_not
g4169 not in1[121] ; in1[121]_not
g4170 not n1759 ; n1759_not
g4171 not n1760 ; n1760_not
g4172 not in1[122] ; in1[122]_not
g4173 not n1762 ; n1762_not
g4174 not n1763 ; n1763_not
g4175 not n1757 ; n1757_not
g4176 not n1764 ; n1764_not
g4177 not n1756 ; n1756_not
g4178 not in0[124] ; in0[124]_not
g4179 not in1[127] ; in1[127]_not
g4180 not in0[126] ; in0[126]_not
g4181 not in0[125] ; in0[125]_not
g4182 not n1769 ; n1769_not
g4183 not n1770 ; n1770_not
g4184 not n1768 ; n1768_not
g4185 not n1767 ; n1767_not
g4186 not n1766 ; n1766_not
g4187 not in1[124] ; in1[124]_not
g4188 not in1[125] ; in1[125]_not
g4189 not n1775 ; n1775_not
g4190 not n1776 ; n1776_not
g4191 not n1777 ; n1777_not
g4192 not in1[126] ; in1[126]_not
g4193 not n1778 ; n1778_not
g4194 not n1779 ; n1779_not
g4195 not n1780 ; n1780_not
g4196 not n1774 ; n1774_not
g4197 not n1781 ; n1781_not
g4198 not n1783 ; n1783_not
g4199 not n1784 ; n1784_not
g4200 not in0[127] ; in0[127]_not
g4201 not n1786 ; n1786_not
g4202 not n1787 ; n1787_not
g4203 not n1788 ; n1788_not
g4204 not n1789 ; n1789_not
g4205 not in2[127] ; in2[127]_not
g4206 not n1791 ; n1791_not
g4207 not n1792 ; n1792_not
g4208 not n1793 ; n1793_not
g4209 not n1794 ; n1794_not
g4210 not n1790 ; n1790_not
g4211 not n1795 ; n1795_not
g4212 not n1798 ; n1798_not
g4213 not n1799 ; n1799_not
g4214 not n1801 ; n1801_not
g4215 not n1802 ; n1802_not
g4216 not n1800 ; n1800_not
g4217 not n1797 ; n1797_not
g4218 not n1804 ; n1804_not
g4219 not n1806 ; n1806_not
g4220 not n1807 ; n1807_not
g4221 not n1809 ; n1809_not
g4222 not n1810 ; n1810_not
g4223 not n1812 ; n1812_not
g4224 not n1813 ; n1813_not
g4225 not n1814 ; n1814_not
g4226 not n1816 ; n1816_not
g4227 not n1817 ; n1817_not
g4228 not n1815 ; n1815_not
g4229 not n1808 ; n1808_not
g4230 not n1811 ; n1811_not
g4231 not n1820 ; n1820_not
g4232 not n1821 ; n1821_not
g4233 not n1822 ; n1822_not
g4234 not n1803 ; n1803_not
g4235 not n1826 ; n1826_not
g4236 not n1827 ; n1827_not
g4237 not n1829 ; n1829_not
g4238 not n1830 ; n1830_not
g4239 not n1828 ; n1828_not
g4240 not n1833 ; n1833_not
g4241 not n1834 ; n1834_not
g4242 not n1836 ; n1836_not
g4243 not n1837 ; n1837_not
g4244 not n1838 ; n1838_not
g4245 not n1840 ; n1840_not
g4246 not n1841 ; n1841_not
g4247 not n1843 ; n1843_not
g4248 not n1844 ; n1844_not
g4249 not n1842 ; n1842_not
g4250 not n1839 ; n1839_not
g4251 not n1846 ; n1846_not
g4252 not n1848 ; n1848_not
g4253 not n1849 ; n1849_not
g4254 not n1851 ; n1851_not
g4255 not n1852 ; n1852_not
g4256 not n1853 ; n1853_not
g4257 not n1855 ; n1855_not
g4258 not n1856 ; n1856_not
g4259 not n1858 ; n1858_not
g4260 not n1859 ; n1859_not
g4261 not n1857 ; n1857_not
g4262 not n1860 ; n1860_not
g4263 not n1863 ; n1863_not
g4264 not n1864 ; n1864_not
g4265 not n1866 ; n1866_not
g4266 not n1867 ; n1867_not
g4267 not n1865 ; n1865_not
g4268 not n1862 ; n1862_not
g4269 not n1869 ; n1869_not
g4270 not n1871 ; n1871_not
g4271 not n1872 ; n1872_not
g4272 not n1874 ; n1874_not
g4273 not n1875 ; n1875_not
g4274 not n1876 ; n1876_not
g4275 not n1878 ; n1878_not
g4276 not n1879 ; n1879_not
g4277 not n1881 ; n1881_not
g4278 not n1882 ; n1882_not
g4279 not n1880 ; n1880_not
g4280 not n1877 ; n1877_not
g4281 not n1873 ; n1873_not
g4282 not n1885 ; n1885_not
g4283 not n1886 ; n1886_not
g4284 not n1887 ; n1887_not
g4285 not n1868 ; n1868_not
g4286 not n1891 ; n1891_not
g4287 not n1892 ; n1892_not
g4288 not n1894 ; n1894_not
g4289 not n1895 ; n1895_not
g4290 not n1893 ; n1893_not
g4291 not n1896 ; n1896_not
g4292 not n1899 ; n1899_not
g4293 not n1900 ; n1900_not
g4294 not n1902 ; n1902_not
g4295 not n1903 ; n1903_not
g4296 not n1901 ; n1901_not
g4297 not n1898 ; n1898_not
g4298 not n1905 ; n1905_not
g4299 not n1907 ; n1907_not
g4300 not n1908 ; n1908_not
g4301 not n1910 ; n1910_not
g4302 not n1911 ; n1911_not
g4303 not n1912 ; n1912_not
g4304 not n1914 ; n1914_not
g4305 not n1915 ; n1915_not
g4306 not n1917 ; n1917_not
g4307 not n1918 ; n1918_not
g4308 not n1916 ; n1916_not
g4309 not n1913 ; n1913_not
g4310 not n1909 ; n1909_not
g4311 not n1921 ; n1921_not
g4312 not n1922 ; n1922_not
g4313 not n1923 ; n1923_not
g4314 not n1904 ; n1904_not
g4315 not n1927 ; n1927_not
g4316 not n1928 ; n1928_not
g4317 not n1930 ; n1930_not
g4318 not n1931 ; n1931_not
g4319 not n1929 ; n1929_not
g4320 not n1934 ; n1934_not
g4321 not n1935 ; n1935_not
g4322 not n1937 ; n1937_not
g4323 not n1938 ; n1938_not
g4324 not n1939 ; n1939_not
g4325 not n1941 ; n1941_not
g4326 not n1942 ; n1942_not
g4327 not n1944 ; n1944_not
g4328 not n1945 ; n1945_not
g4329 not n1943 ; n1943_not
g4330 not n1940 ; n1940_not
g4331 not n1947 ; n1947_not
g4332 not n1949 ; n1949_not
g4333 not n1950 ; n1950_not
g4334 not n1952 ; n1952_not
g4335 not n1953 ; n1953_not
g4336 not n1954 ; n1954_not
g4337 not n1956 ; n1956_not
g4338 not n1957 ; n1957_not
g4339 not n1959 ; n1959_not
g4340 not n1960 ; n1960_not
g4341 not n1958 ; n1958_not
g4342 not n1961 ; n1961_not
g4343 not n1964 ; n1964_not
g4344 not n1965 ; n1965_not
g4345 not n1967 ; n1967_not
g4346 not n1968 ; n1968_not
g4347 not n1966 ; n1966_not
g4348 not n1963 ; n1963_not
g4349 not n1970 ; n1970_not
g4350 not n1972 ; n1972_not
g4351 not n1973 ; n1973_not
g4352 not n1975 ; n1975_not
g4353 not n1976 ; n1976_not
g4354 not n1977 ; n1977_not
g4355 not n1979 ; n1979_not
g4356 not n1980 ; n1980_not
g4357 not n1982 ; n1982_not
g4358 not n1983 ; n1983_not
g4359 not n1981 ; n1981_not
g4360 not n1978 ; n1978_not
g4361 not n1974 ; n1974_not
g4362 not n1986 ; n1986_not
g4363 not n1987 ; n1987_not
g4364 not n1988 ; n1988_not
g4365 not n1969 ; n1969_not
g4366 not n1992 ; n1992_not
g4367 not n1993 ; n1993_not
g4368 not n1995 ; n1995_not
g4369 not n1996 ; n1996_not
g4370 not n1994 ; n1994_not
g4371 not n1997 ; n1997_not
g4372 not n2000 ; n2000_not
g4373 not n2001 ; n2001_not
g4374 not n2003 ; n2003_not
g4375 not n2004 ; n2004_not
g4376 not n2002 ; n2002_not
g4377 not n1999 ; n1999_not
g4378 not n2006 ; n2006_not
g4379 not n2008 ; n2008_not
g4380 not n2009 ; n2009_not
g4381 not n2011 ; n2011_not
g4382 not n2012 ; n2012_not
g4383 not n2013 ; n2013_not
g4384 not n2015 ; n2015_not
g4385 not n2016 ; n2016_not
g4386 not n2018 ; n2018_not
g4387 not n2019 ; n2019_not
g4388 not n2017 ; n2017_not
g4389 not n2014 ; n2014_not
g4390 not n2010 ; n2010_not
g4391 not n2022 ; n2022_not
g4392 not n2023 ; n2023_not
g4393 not n2024 ; n2024_not
g4394 not n2005 ; n2005_not
g4395 not n2028 ; n2028_not
g4396 not n2029 ; n2029_not
g4397 not n2031 ; n2031_not
g4398 not n2032 ; n2032_not
g4399 not n2030 ; n2030_not
g4400 not n2035 ; n2035_not
g4401 not n2036 ; n2036_not
g4402 not n2038 ; n2038_not
g4403 not n2039 ; n2039_not
g4404 not n2040 ; n2040_not
g4405 not n2042 ; n2042_not
g4406 not n2043 ; n2043_not
g4407 not n2045 ; n2045_not
g4408 not n2046 ; n2046_not
g4409 not n2044 ; n2044_not
g4410 not n2041 ; n2041_not
g4411 not n2048 ; n2048_not
g4412 not n2050 ; n2050_not
g4413 not n2051 ; n2051_not
g4414 not n2053 ; n2053_not
g4415 not n2054 ; n2054_not
g4416 not n2055 ; n2055_not
g4417 not n2057 ; n2057_not
g4418 not n2058 ; n2058_not
g4419 not n2060 ; n2060_not
g4420 not n2061 ; n2061_not
g4421 not n2059 ; n2059_not
g4422 not n2062 ; n2062_not
g4423 not n2065 ; n2065_not
g4424 not n2066 ; n2066_not
g4425 not n2068 ; n2068_not
g4426 not n2069 ; n2069_not
g4427 not n2067 ; n2067_not
g4428 not n2064 ; n2064_not
g4429 not n2071 ; n2071_not
g4430 not n2073 ; n2073_not
g4431 not n2074 ; n2074_not
g4432 not n2076 ; n2076_not
g4433 not n2077 ; n2077_not
g4434 not n2078 ; n2078_not
g4435 not n2080 ; n2080_not
g4436 not n2081 ; n2081_not
g4437 not n2083 ; n2083_not
g4438 not n2084 ; n2084_not
g4439 not n2082 ; n2082_not
g4440 not n2079 ; n2079_not
g4441 not n2075 ; n2075_not
g4442 not n2087 ; n2087_not
g4443 not n2088 ; n2088_not
g4444 not n2089 ; n2089_not
g4445 not n2070 ; n2070_not
g4446 not n2093 ; n2093_not
g4447 not n2094 ; n2094_not
g4448 not n2096 ; n2096_not
g4449 not n2097 ; n2097_not
g4450 not n2095 ; n2095_not
g4451 not n2098 ; n2098_not
g4452 not n2101 ; n2101_not
g4453 not n2102 ; n2102_not
g4454 not n2104 ; n2104_not
g4455 not n2105 ; n2105_not
g4456 not n2103 ; n2103_not
g4457 not n2100 ; n2100_not
g4458 not n2107 ; n2107_not
g4459 not n2109 ; n2109_not
g4460 not n2110 ; n2110_not
g4461 not n2112 ; n2112_not
g4462 not n2113 ; n2113_not
g4463 not n2114 ; n2114_not
g4464 not n2116 ; n2116_not
g4465 not n2117 ; n2117_not
g4466 not n2119 ; n2119_not
g4467 not n2120 ; n2120_not
g4468 not n2118 ; n2118_not
g4469 not n2115 ; n2115_not
g4470 not n2111 ; n2111_not
g4471 not n2123 ; n2123_not
g4472 not n2124 ; n2124_not
g4473 not n2125 ; n2125_not
g4474 not n2106 ; n2106_not
g4475 not n2129 ; n2129_not
g4476 not n2130 ; n2130_not
g4477 not n2132 ; n2132_not
g4478 not n2133 ; n2133_not
g4479 not n2134 ; n2134_not
g4480 not n2136 ; n2136_not
g4481 not n2137 ; n2137_not
g4482 not n2139 ; n2139_not
g4483 not n2140 ; n2140_not
g4484 not n2138 ; n2138_not
g4485 not n2135 ; n2135_not
g4486 not n2142 ; n2142_not
g4487 not n2144 ; n2144_not
g4488 not n2145 ; n2145_not
g4489 not n2147 ; n2147_not
g4490 not n2148 ; n2148_not
g4491 not n2146 ; n2146_not
g4492 not n2151 ; n2151_not
g4493 not n2152 ; n2152_not
g4494 not n2154 ; n2154_not
g4495 not n2155 ; n2155_not
g4496 not n2156 ; n2156_not
g4497 not n2158 ; n2158_not
g4498 not n2159 ; n2159_not
g4499 not n2161 ; n2161_not
g4500 not n2162 ; n2162_not
g4501 not n2160 ; n2160_not
g4502 not n2163 ; n2163_not
g4503 not n2166 ; n2166_not
g4504 not n2167 ; n2167_not
g4505 not n2169 ; n2169_not
g4506 not n2170 ; n2170_not
g4507 not n2168 ; n2168_not
g4508 not n2165 ; n2165_not
g4509 not n2172 ; n2172_not
g4510 not n2174 ; n2174_not
g4511 not n2175 ; n2175_not
g4512 not n2177 ; n2177_not
g4513 not n2178 ; n2178_not
g4514 not n2179 ; n2179_not
g4515 not n2181 ; n2181_not
g4516 not n2182 ; n2182_not
g4517 not n2184 ; n2184_not
g4518 not n2185 ; n2185_not
g4519 not n2186 ; n2186_not
g4520 not n2180 ; n2180_not
g4521 not n2187 ; n2187_not
g4522 not n2190 ; n2190_not
g4523 not n2191 ; n2191_not
g4524 not n2193 ; n2193_not
g4525 not n2194 ; n2194_not
g4526 not n2192 ; n2192_not
g4527 not n2195 ; n2195_not
g4528 not n2198 ; n2198_not
g4529 not n2199 ; n2199_not
g4530 not n2201 ; n2201_not
g4531 not n2202 ; n2202_not
g4532 not n2203 ; n2203_not
g4533 not n2197 ; n2197_not
g4534 not n2204 ; n2204_not
g4535 not n2206 ; n2206_not
g4536 not n2207 ; n2207_not
g4537 not n2209 ; n2209_not
g4538 not n2210 ; n2210_not
g4539 not n2211 ; n2211_not
g4540 not n2213 ; n2213_not
g4541 not n2214 ; n2214_not
g4542 not n2216 ; n2216_not
g4543 not n2217 ; n2217_not
g4544 not n2215 ; n2215_not
g4545 not n2212 ; n2212_not
g4546 not n2208 ; n2208_not
g4547 not n2220 ; n2220_not
g4548 not n2221 ; n2221_not
g4549 not n2200 ; n2200_not
g4550 not n2223 ; n2223_not
g4551 not n2224 ; n2224_not
g4552 not n2196 ; n2196_not
g4553 not n2225 ; n2225_not
g4554 not n2226 ; n2226_not
g4555 not n2176 ; n2176_not
g4556 not n2183 ; n2183_not
g4557 not n2229 ; n2229_not
g4558 not n2230 ; n2230_not
g4559 not n2231 ; n2231_not
g4560 not n2171 ; n2171_not
g4561 not n2235 ; n2235_not
g4562 not n2236 ; n2236_not
g4563 not n2238 ; n2238_not
g4564 not n2239 ; n2239_not
g4565 not n2237 ; n2237_not
g4566 not n2240 ; n2240_not
g4567 not n2243 ; n2243_not
g4568 not n2244 ; n2244_not
g4569 not n2246 ; n2246_not
g4570 not n2247 ; n2247_not
g4571 not n2245 ; n2245_not
g4572 not n2242 ; n2242_not
g4573 not n2249 ; n2249_not
g4574 not n2251 ; n2251_not
g4575 not n2252 ; n2252_not
g4576 not n2254 ; n2254_not
g4577 not n2255 ; n2255_not
g4578 not n2256 ; n2256_not
g4579 not n2258 ; n2258_not
g4580 not n2259 ; n2259_not
g4581 not n2261 ; n2261_not
g4582 not n2262 ; n2262_not
g4583 not n2263 ; n2263_not
g4584 not n2257 ; n2257_not
g4585 not n2264 ; n2264_not
g4586 not n2267 ; n2267_not
g4587 not n2268 ; n2268_not
g4588 not n2270 ; n2270_not
g4589 not n2271 ; n2271_not
g4590 not n2269 ; n2269_not
g4591 not n2272 ; n2272_not
g4592 not n2275 ; n2275_not
g4593 not n2276 ; n2276_not
g4594 not n2278 ; n2278_not
g4595 not n2279 ; n2279_not
g4596 not n2280 ; n2280_not
g4597 not n2274 ; n2274_not
g4598 not n2281 ; n2281_not
g4599 not n2283 ; n2283_not
g4600 not n2284 ; n2284_not
g4601 not n2286 ; n2286_not
g4602 not n2287 ; n2287_not
g4603 not n2288 ; n2288_not
g4604 not n2290 ; n2290_not
g4605 not n2291 ; n2291_not
g4606 not n2293 ; n2293_not
g4607 not n2294 ; n2294_not
g4608 not n2292 ; n2292_not
g4609 not n2289 ; n2289_not
g4610 not n2285 ; n2285_not
g4611 not n2297 ; n2297_not
g4612 not n2298 ; n2298_not
g4613 not n2277 ; n2277_not
g4614 not n2300 ; n2300_not
g4615 not n2301 ; n2301_not
g4616 not n2273 ; n2273_not
g4617 not n2302 ; n2302_not
g4618 not n2303 ; n2303_not
g4619 not n2253 ; n2253_not
g4620 not n2260 ; n2260_not
g4621 not n2306 ; n2306_not
g4622 not n2307 ; n2307_not
g4623 not n2308 ; n2308_not
g4624 not n2248 ; n2248_not
g4625 not n2312 ; n2312_not
g4626 not n2313 ; n2313_not
g4627 not n2315 ; n2315_not
g4628 not n2316 ; n2316_not
g4629 not n2314 ; n2314_not
g4630 not n2319 ; n2319_not
g4631 not n2320 ; n2320_not
g4632 not n2322 ; n2322_not
g4633 not n2323 ; n2323_not
g4634 not n2324 ; n2324_not
g4635 not n2326 ; n2326_not
g4636 not n2327 ; n2327_not
g4637 not n2329 ; n2329_not
g4638 not n2330 ; n2330_not
g4639 not n2331 ; n2331_not
g4640 not n2333 ; n2333_not
g4641 not n2334 ; n2334_not
g4642 not n2336 ; n2336_not
g4643 not n2337 ; n2337_not
g4644 not n2338 ; n2338_not
g4645 not n2340 ; n2340_not
g4646 not n2341 ; n2341_not
g4647 not n2343 ; n2343_not
g4648 not n2344 ; n2344_not
g4649 not n2345 ; n2345_not
g4650 not n2347 ; n2347_not
g4651 not n2348 ; n2348_not
g4652 not n2350 ; n2350_not
g4653 not n2351 ; n2351_not
g4654 not n2352 ; n2352_not
g4655 not n2354 ; n2354_not
g4656 not n2355 ; n2355_not
g4657 not n2357 ; n2357_not
g4658 not n2358 ; n2358_not
g4659 not n2359 ; n2359_not
g4660 not n2361 ; n2361_not
g4661 not n2362 ; n2362_not
g4662 not n2364 ; n2364_not
g4663 not n2365 ; n2365_not
g4664 not n2367 ; n2367_not
g4665 not n2368 ; n2368_not
g4666 not n2370 ; n2370_not
g4667 not n2371 ; n2371_not
g4668 not n2372 ; n2372_not
g4669 not n2374 ; n2374_not
g4670 not n2375 ; n2375_not
g4671 not n2377 ; n2377_not
g4672 not n2378 ; n2378_not
g4673 not n2379 ; n2379_not
g4674 not n2381 ; n2381_not
g4675 not n2382 ; n2382_not
g4676 not n2384 ; n2384_not
g4677 not n2385 ; n2385_not
g4678 not n2386 ; n2386_not
g4679 not n2388 ; n2388_not
g4680 not n2389 ; n2389_not
g4681 not n2391 ; n2391_not
g4682 not n2392 ; n2392_not
g4683 not n2393 ; n2393_not
g4684 not n2395 ; n2395_not
g4685 not n2396 ; n2396_not
g4686 not n2398 ; n2398_not
g4687 not n2399 ; n2399_not
g4688 not n2400 ; n2400_not
g4689 not n2402 ; n2402_not
g4690 not n2403 ; n2403_not
g4691 not n2405 ; n2405_not
g4692 not n2406 ; n2406_not
g4693 not n2407 ; n2407_not
g4694 not n2409 ; n2409_not
g4695 not n2410 ; n2410_not
g4696 not n2412 ; n2412_not
g4697 not n2413 ; n2413_not
g4698 not n2415 ; n2415_not
g4699 not n2416 ; n2416_not
g4700 not n2418 ; n2418_not
g4701 not n2419 ; n2419_not
g4702 not n2420 ; n2420_not
g4703 not n2422 ; n2422_not
g4704 not n2423 ; n2423_not
g4705 not n2425 ; n2425_not
g4706 not n2426 ; n2426_not
g4707 not n2427 ; n2427_not
g4708 not n2429 ; n2429_not
g4709 not n2430 ; n2430_not
g4710 not n2432 ; n2432_not
g4711 not n2433 ; n2433_not
g4712 not n2434 ; n2434_not
g4713 not n2436 ; n2436_not
g4714 not n2437 ; n2437_not
g4715 not n2439 ; n2439_not
g4716 not n2440 ; n2440_not
g4717 not n2441 ; n2441_not
g4718 not n2443 ; n2443_not
g4719 not n2444 ; n2444_not
g4720 not n2446 ; n2446_not
g4721 not n2447 ; n2447_not
g4722 not n2448 ; n2448_not
g4723 not n2450 ; n2450_not
g4724 not n2451 ; n2451_not
g4725 not n2453 ; n2453_not
g4726 not n2454 ; n2454_not
g4727 not n2455 ; n2455_not
g4728 not n2457 ; n2457_not
g4729 not n2458 ; n2458_not
g4730 not n2460 ; n2460_not
g4731 not n2461 ; n2461_not
g4732 not n2463 ; n2463_not
g4733 not n2464 ; n2464_not
g4734 not n2466 ; n2466_not
g4735 not n2467 ; n2467_not
g4736 not n2468 ; n2468_not
g4737 not n2470 ; n2470_not
g4738 not n2471 ; n2471_not
g4739 not n2473 ; n2473_not
g4740 not n2474 ; n2474_not
g4741 not n2476 ; n2476_not
g4742 not n2477 ; n2477_not
g4743 not n2479 ; n2479_not
g4744 not n2480 ; n2480_not
g4745 not n2482 ; n2482_not
g4746 not n2483 ; n2483_not
g4747 not n2485 ; n2485_not
g4748 not n2486 ; n2486_not
g4749 not n2488 ; n2488_not
g4750 not n2489 ; n2489_not
g4751 not n2491 ; n2491_not
g4752 not n2492 ; n2492_not
g4753 not n2493 ; n2493_not
g4754 not n2495 ; n2495_not
g4755 not n2496 ; n2496_not
g4756 not n2498 ; n2498_not
g4757 not n2499 ; n2499_not
g4758 not n2501 ; n2501_not
g4759 not n2502 ; n2502_not
g4760 not n2500 ; n2500_not
g4761 not n2506 ; n2506_not
g4762 not n2507 ; n2507_not
g4763 not n2505 ; n2505_not
g4764 not n2510 ; n2510_not
g4765 not n2511 ; n2511_not
g4766 not n2513 ; n2513_not
g4767 not n2514 ; n2514_not
g4768 not n2515 ; n2515_not
g4769 not n2497 ; n2497_not
g4770 not n2504 ; n2504_not
g4771 not n2516 ; n2516_not
g4772 not n2517 ; n2517_not
g4773 not n2509 ; n2509_not
g4774 not n2512 ; n2512_not
g4775 not n2519 ; n2519_not
g4776 not n2520 ; n2520_not
g4777 not n2494 ; n2494_not
g4778 not n2521 ; n2521_not
g4779 not n2490 ; n2490_not
g4780 not n2522 ; n2522_not
g4781 not n2523 ; n2523_not
g4782 not n2525 ; n2525_not
g4783 not n2487 ; n2487_not
g4784 not n2524 ; n2524_not
g4785 not n2526 ; n2526_not
g4786 not n2527 ; n2527_not
g4787 not n2529 ; n2529_not
g4788 not n2481 ; n2481_not
g4789 not n2528 ; n2528_not
g4790 not n2530 ; n2530_not
g4791 not n2531 ; n2531_not
g4792 not n2533 ; n2533_not
g4793 not n2475 ; n2475_not
g4794 not n2532 ; n2532_not
g4795 not n2534 ; n2534_not
g4796 not n2535 ; n2535_not
g4797 not n2469 ; n2469_not
g4798 not n2536 ; n2536_not
g4799 not n2465 ; n2465_not
g4800 not n2537 ; n2537_not
g4801 not n2538 ; n2538_not
g4802 not n2540 ; n2540_not
g4803 not n2541 ; n2541_not
g4804 not n2543 ; n2543_not
g4805 not n2539 ; n2539_not
g4806 not n2542 ; n2542_not
g4807 not n2544 ; n2544_not
g4808 not n2545 ; n2545_not
g4809 not n2547 ; n2547_not
g4810 not n2548 ; n2548_not
g4811 not n2550 ; n2550_not
g4812 not n2546 ; n2546_not
g4813 not n2549 ; n2549_not
g4814 not n2551 ; n2551_not
g4815 not n2552 ; n2552_not
g4816 not n2456 ; n2456_not
g4817 not n2553 ; n2553_not
g4818 not n2452 ; n2452_not
g4819 not n2554 ; n2554_not
g4820 not n2555 ; n2555_not
g4821 not n2449 ; n2449_not
g4822 not n2556 ; n2556_not
g4823 not n2445 ; n2445_not
g4824 not n2557 ; n2557_not
g4825 not n2558 ; n2558_not
g4826 not n2442 ; n2442_not
g4827 not n2559 ; n2559_not
g4828 not n2438 ; n2438_not
g4829 not n2560 ; n2560_not
g4830 not n2561 ; n2561_not
g4831 not n2435 ; n2435_not
g4832 not n2562 ; n2562_not
g4833 not n2431 ; n2431_not
g4834 not n2563 ; n2563_not
g4835 not n2564 ; n2564_not
g4836 not n2428 ; n2428_not
g4837 not n2565 ; n2565_not
g4838 not n2424 ; n2424_not
g4839 not n2566 ; n2566_not
g4840 not n2567 ; n2567_not
g4841 not n2421 ; n2421_not
g4842 not n2568 ; n2568_not
g4843 not n2417 ; n2417_not
g4844 not n2569 ; n2569_not
g4845 not n2570 ; n2570_not
g4846 not n2572 ; n2572_not
g4847 not n2573 ; n2573_not
g4848 not n2575 ; n2575_not
g4849 not n2571 ; n2571_not
g4850 not n2574 ; n2574_not
g4851 not n2576 ; n2576_not
g4852 not n2577 ; n2577_not
g4853 not n2579 ; n2579_not
g4854 not n2580 ; n2580_not
g4855 not n2582 ; n2582_not
g4856 not n2578 ; n2578_not
g4857 not n2581 ; n2581_not
g4858 not n2583 ; n2583_not
g4859 not n2584 ; n2584_not
g4860 not n2408 ; n2408_not
g4861 not n2585 ; n2585_not
g4862 not n2404 ; n2404_not
g4863 not n2586 ; n2586_not
g4864 not n2587 ; n2587_not
g4865 not n2401 ; n2401_not
g4866 not n2588 ; n2588_not
g4867 not n2397 ; n2397_not
g4868 not n2589 ; n2589_not
g4869 not n2590 ; n2590_not
g4870 not n2394 ; n2394_not
g4871 not n2591 ; n2591_not
g4872 not n2390 ; n2390_not
g4873 not n2592 ; n2592_not
g4874 not n2593 ; n2593_not
g4875 not n2387 ; n2387_not
g4876 not n2594 ; n2594_not
g4877 not n2383 ; n2383_not
g4878 not n2595 ; n2595_not
g4879 not n2596 ; n2596_not
g4880 not n2380 ; n2380_not
g4881 not n2597 ; n2597_not
g4882 not n2376 ; n2376_not
g4883 not n2598 ; n2598_not
g4884 not n2599 ; n2599_not
g4885 not n2373 ; n2373_not
g4886 not n2600 ; n2600_not
g4887 not n2369 ; n2369_not
g4888 not n2601 ; n2601_not
g4889 not n2602 ; n2602_not
g4890 not n2604 ; n2604_not
g4891 not n2605 ; n2605_not
g4892 not n2607 ; n2607_not
g4893 not n2603 ; n2603_not
g4894 not n2606 ; n2606_not
g4895 not n2608 ; n2608_not
g4896 not n2609 ; n2609_not
g4897 not n2611 ; n2611_not
g4898 not n2612 ; n2612_not
g4899 not n2614 ; n2614_not
g4900 not n2610 ; n2610_not
g4901 not n2613 ; n2613_not
g4902 not n2615 ; n2615_not
g4903 not n2616 ; n2616_not
g4904 not n2360 ; n2360_not
g4905 not n2617 ; n2617_not
g4906 not n2356 ; n2356_not
g4907 not n2618 ; n2618_not
g4908 not n2619 ; n2619_not
g4909 not n2353 ; n2353_not
g4910 not n2620 ; n2620_not
g4911 not n2349 ; n2349_not
g4912 not n2621 ; n2621_not
g4913 not n2622 ; n2622_not
g4914 not n2346 ; n2346_not
g4915 not n2623 ; n2623_not
g4916 not n2342 ; n2342_not
g4917 not n2624 ; n2624_not
g4918 not n2625 ; n2625_not
g4919 not n2339 ; n2339_not
g4920 not n2626 ; n2626_not
g4921 not n2335 ; n2335_not
g4922 not n2627 ; n2627_not
g4923 not n2628 ; n2628_not
g4924 not n2332 ; n2332_not
g4925 not n2629 ; n2629_not
g4926 not n2328 ; n2328_not
g4927 not n2630 ; n2630_not
g4928 not n2631 ; n2631_not
g4929 not n2325 ; n2325_not
g4930 not n2632 ; n2632_not
g4931 not n2321 ; n2321_not
g4932 not n2633 ; n2633_not
g4933 not n2634 ; n2634_not
g4934 not n2636 ; n2636_not
g4935 not n2637 ; n2637_not
g4936 not n2639 ; n2639_not
g4937 not n2640 ; n2640_not
g4938 not n2641 ; n2641_not
g4939 not n2643 ; n2643_not
g4940 not n2644 ; n2644_not
g4941 not n2646 ; n2646_not
g4942 not n2647 ; n2647_not
g4943 not n2645 ; n2645_not
g4944 not n2642 ; n2642_not
g4945 not n2649 ; n2649_not
g4946 not n2651 ; n2651_not
g4947 not n2652 ; n2652_not
g4948 not n2654 ; n2654_not
g4949 not n2655 ; n2655_not
g4950 not n2656 ; n2656_not
g4951 not n2658 ; n2658_not
g4952 not n2659 ; n2659_not
g4953 not n2661 ; n2661_not
g4954 not n2662 ; n2662_not
g4955 not n2663 ; n2663_not
g4956 not n2657 ; n2657_not
g4957 not n2664 ; n2664_not
g4958 not n2667 ; n2667_not
g4959 not n2668 ; n2668_not
g4960 not n2670 ; n2670_not
g4961 not n2671 ; n2671_not
g4962 not n2672 ; n2672_not
g4963 not n2674 ; n2674_not
g4964 not n2675 ; n2675_not
g4965 not n2677 ; n2677_not
g4966 not n2678 ; n2678_not
g4967 not n2679 ; n2679_not
g4968 not n2681 ; n2681_not
g4969 not n2682 ; n2682_not
g4970 not n2684 ; n2684_not
g4971 not n2685 ; n2685_not
g4972 not n2683 ; n2683_not
g4973 not n2680 ; n2680_not
g4974 not n2687 ; n2687_not
g4975 not n2673 ; n2673_not
g4976 not n2635 ; n2635_not
g4977 not n2318 ; n2318_not
g4978 not n2638 ; n2638_not
g4979 not n2653 ; n2653_not
g4980 not n2660 ; n2660_not
g4981 not n2695 ; n2695_not
g4982 not n2696 ; n2696_not
g4983 not n2697 ; n2697_not
g4984 not n2648 ; n2648_not
g4985 not n2676 ; n2676_not
g4986 not n2686 ; n2686_not
g4987 not n2317 ; n2317_not
g4988 not n2669 ; n2669_not
g4989 not n2704 ; n2704_not
g4990 not n2705 ; n2705_not
g4991 not n2706 ; n2706_not
g4992 not n2703 ; n2703_not
g4993 not n2707 ; n2707_not
g4994 not n2701 ; n2701_not
g4995 not n2709 ; n2709_not
g4996 not n2700 ; n2700_not
g4997 not n2710 ; n2710_not
g4998 not n2698 ; n2698_not
g4999 not n2693 ; n2693_not
g5000 not n2692 ; n2692_not
g5001 not n2295 ; n2295_not
g5002 not n2715 ; n2715_not
g5003 not n2714 ; n2714_not
g5004 not n2311 ; n2311_not
g5005 not n2719 ; n2719_not
g5006 not n2309 ; n2309_not
g5007 not n2304 ; n2304_not
g5008 not n2241 ; n2241_not
g5009 not n2724 ; n2724_not
g5010 not n2725 ; n2725_not
g5011 not n2727 ; n2727_not
g5012 not n2728 ; n2728_not
g5013 not n2726 ; n2726_not
g5014 not n2731 ; n2731_not
g5015 not n2732 ; n2732_not
g5016 not n2734 ; n2734_not
g5017 not n2735 ; n2735_not
g5018 not n2736 ; n2736_not
g5019 not n2738 ; n2738_not
g5020 not n2739 ; n2739_not
g5021 not n2741 ; n2741_not
g5022 not n2742 ; n2742_not
g5023 not n2740 ; n2740_not
g5024 not n2737 ; n2737_not
g5025 not n2744 ; n2744_not
g5026 not n2746 ; n2746_not
g5027 not n2747 ; n2747_not
g5028 not n2749 ; n2749_not
g5029 not n2750 ; n2750_not
g5030 not n2751 ; n2751_not
g5031 not n2753 ; n2753_not
g5032 not n2754 ; n2754_not
g5033 not n2756 ; n2756_not
g5034 not n2757 ; n2757_not
g5035 not n2755 ; n2755_not
g5036 not n2752 ; n2752_not
g5037 not n2759 ; n2759_not
g5038 not n2762 ; n2762_not
g5039 not n2763 ; n2763_not
g5040 not n2765 ; n2765_not
g5041 not n2766 ; n2766_not
g5042 not n2767 ; n2767_not
g5043 not n2769 ; n2769_not
g5044 not n2770 ; n2770_not
g5045 not n2772 ; n2772_not
g5046 not n2773 ; n2773_not
g5047 not n2774 ; n2774_not
g5048 not n2776 ; n2776_not
g5049 not n2777 ; n2777_not
g5050 not n2779 ; n2779_not
g5051 not n2780 ; n2780_not
g5052 not n2778 ; n2778_not
g5053 not n2775 ; n2775_not
g5054 not n2782 ; n2782_not
g5055 not n2768 ; n2768_not
g5056 not n2730 ; n2730_not
g5057 not n2723 ; n2723_not
g5058 not n2733 ; n2733_not
g5059 not n2771 ; n2771_not
g5060 not n2781 ; n2781_not
g5061 not n2729 ; n2729_not
g5062 not n2764 ; n2764_not
g5063 not n2792 ; n2792_not
g5064 not n2793 ; n2793_not
g5065 not n2794 ; n2794_not
g5066 not n2791 ; n2791_not
g5067 not n2795 ; n2795_not
g5068 not n2789 ; n2789_not
g5069 not n2797 ; n2797_not
g5070 not n2758 ; n2758_not
g5071 not n2748 ; n2748_not
g5072 not n2800 ; n2800_not
g5073 not n2801 ; n2801_not
g5074 not n2743 ; n2743_not
g5075 not n2803 ; n2803_not
g5076 not n2804 ; n2804_not
g5077 not n2798 ; n2798_not
g5078 not n2805 ; n2805_not
g5079 not n2788 ; n2788_not
g5080 not n2787 ; n2787_not
g5081 not n2218 ; n2218_not
g5082 not n2809 ; n2809_not
g5083 not n2808 ; n2808_not
g5084 not n2234 ; n2234_not
g5085 not n2813 ; n2813_not
g5086 not n2232 ; n2232_not
g5087 not n2227 ; n2227_not
g5088 not n2164 ; n2164_not
g5089 not n2157 ; n2157_not
g5090 not n2817 ; n2817_not
g5091 not n2150 ; n2150_not
g5092 not n2131 ; n2131_not
g5093 not n2149 ; n2149_not
g5094 not n2153 ; n2153_not
g5095 not n2823 ; n2823_not
g5096 not n2824 ; n2824_not
g5097 not n2141 ; n2141_not
g5098 not n2826 ; n2826_not
g5099 not n2827 ; n2827_not
g5100 not n2821 ; n2821_not
g5101 not n2828 ; n2828_not
g5102 not n2820 ; n2820_not
g5103 not n2121 ; n2121_not
g5104 not n2831 ; n2831_not
g5105 not n2830 ; n2830_not
g5106 not n2128 ; n2128_not
g5107 not n2834 ; n2834_not
g5108 not n2126 ; n2126_not
g5109 not n2099 ; n2099_not
g5110 not n2838 ; n2838_not
g5111 not n2839 ; n2839_not
g5112 not n2841 ; n2841_not
g5113 not n2842 ; n2842_not
g5114 not n2843 ; n2843_not
g5115 not n2845 ; n2845_not
g5116 not n2846 ; n2846_not
g5117 not n2848 ; n2848_not
g5118 not n2849 ; n2849_not
g5119 not n2847 ; n2847_not
g5120 not n2844 ; n2844_not
g5121 not n2851 ; n2851_not
g5122 not n2853 ; n2853_not
g5123 not n2854 ; n2854_not
g5124 not n2856 ; n2856_not
g5125 not n2857 ; n2857_not
g5126 not n2858 ; n2858_not
g5127 not n2860 ; n2860_not
g5128 not n2861 ; n2861_not
g5129 not n2863 ; n2863_not
g5130 not n2864 ; n2864_not
g5131 not n2862 ; n2862_not
g5132 not n2859 ; n2859_not
g5133 not n2866 ; n2866_not
g5134 not n2837 ; n2837_not
g5135 not n2840 ; n2840_not
g5136 not n2865 ; n2865_not
g5137 not n2855 ; n2855_not
g5138 not n2872 ; n2872_not
g5139 not n2873 ; n2873_not
g5140 not n2850 ; n2850_not
g5141 not n2875 ; n2875_not
g5142 not n2876 ; n2876_not
g5143 not n2870 ; n2870_not
g5144 not n2877 ; n2877_not
g5145 not n2869 ; n2869_not
g5146 not n2085 ; n2085_not
g5147 not n2880 ; n2880_not
g5148 not n2879 ; n2879_not
g5149 not n2092 ; n2092_not
g5150 not n2883 ; n2883_not
g5151 not n2090 ; n2090_not
g5152 not n2063 ; n2063_not
g5153 not n2056 ; n2056_not
g5154 not n2886 ; n2886_not
g5155 not n2034 ; n2034_not
g5156 not n2037 ; n2037_not
g5157 not n2033 ; n2033_not
g5158 not n2052 ; n2052_not
g5159 not n2892 ; n2892_not
g5160 not n2893 ; n2893_not
g5161 not n2047 ; n2047_not
g5162 not n2895 ; n2895_not
g5163 not n2896 ; n2896_not
g5164 not n2890 ; n2890_not
g5165 not n2897 ; n2897_not
g5166 not n2889 ; n2889_not
g5167 not n2020 ; n2020_not
g5168 not n2900 ; n2900_not
g5169 not n2899 ; n2899_not
g5170 not n2027 ; n2027_not
g5171 not n2903 ; n2903_not
g5172 not n2025 ; n2025_not
g5173 not n1998 ; n1998_not
g5174 not n2907 ; n2907_not
g5175 not n2908 ; n2908_not
g5176 not n2910 ; n2910_not
g5177 not n2911 ; n2911_not
g5178 not n2912 ; n2912_not
g5179 not n2914 ; n2914_not
g5180 not n2915 ; n2915_not
g5181 not n2917 ; n2917_not
g5182 not n2918 ; n2918_not
g5183 not n2916 ; n2916_not
g5184 not n2913 ; n2913_not
g5185 not n2920 ; n2920_not
g5186 not n2922 ; n2922_not
g5187 not n2923 ; n2923_not
g5188 not n2925 ; n2925_not
g5189 not n2926 ; n2926_not
g5190 not n2927 ; n2927_not
g5191 not n2929 ; n2929_not
g5192 not n2930 ; n2930_not
g5193 not n2932 ; n2932_not
g5194 not n2933 ; n2933_not
g5195 not n2931 ; n2931_not
g5196 not n2928 ; n2928_not
g5197 not n2935 ; n2935_not
g5198 not n2906 ; n2906_not
g5199 not n2909 ; n2909_not
g5200 not n2934 ; n2934_not
g5201 not n2924 ; n2924_not
g5202 not n2941 ; n2941_not
g5203 not n2942 ; n2942_not
g5204 not n2919 ; n2919_not
g5205 not n2944 ; n2944_not
g5206 not n2945 ; n2945_not
g5207 not n2939 ; n2939_not
g5208 not n2946 ; n2946_not
g5209 not n2938 ; n2938_not
g5210 not n1984 ; n1984_not
g5211 not n2949 ; n2949_not
g5212 not n2948 ; n2948_not
g5213 not n1991 ; n1991_not
g5214 not n2952 ; n2952_not
g5215 not n1989 ; n1989_not
g5216 not n1962 ; n1962_not
g5217 not n1955 ; n1955_not
g5218 not n2955 ; n2955_not
g5219 not n1933 ; n1933_not
g5220 not n1936 ; n1936_not
g5221 not n1932 ; n1932_not
g5222 not n1951 ; n1951_not
g5223 not n2961 ; n2961_not
g5224 not n2962 ; n2962_not
g5225 not n1946 ; n1946_not
g5226 not n2964 ; n2964_not
g5227 not n2965 ; n2965_not
g5228 not n2959 ; n2959_not
g5229 not n2966 ; n2966_not
g5230 not n2958 ; n2958_not
g5231 not n1919 ; n1919_not
g5232 not n2969 ; n2969_not
g5233 not n2968 ; n2968_not
g5234 not n1926 ; n1926_not
g5235 not n2972 ; n2972_not
g5236 not n1924 ; n1924_not
g5237 not n1897 ; n1897_not
g5238 not n2976 ; n2976_not
g5239 not n2977 ; n2977_not
g5240 not n2979 ; n2979_not
g5241 not n2980 ; n2980_not
g5242 not n2981 ; n2981_not
g5243 not n2983 ; n2983_not
g5244 not n2984 ; n2984_not
g5245 not n2986 ; n2986_not
g5246 not n2987 ; n2987_not
g5247 not n2985 ; n2985_not
g5248 not n2982 ; n2982_not
g5249 not n2989 ; n2989_not
g5250 not n2991 ; n2991_not
g5251 not n2992 ; n2992_not
g5252 not n2994 ; n2994_not
g5253 not n2995 ; n2995_not
g5254 not n2996 ; n2996_not
g5255 not n2998 ; n2998_not
g5256 not n2999 ; n2999_not
g5257 not n3001 ; n3001_not
g5258 not n3002 ; n3002_not
g5259 not n3000 ; n3000_not
g5260 not n2997 ; n2997_not
g5261 not n3004 ; n3004_not
g5262 not n2975 ; n2975_not
g5263 not n2978 ; n2978_not
g5264 not n3003 ; n3003_not
g5265 not n2993 ; n2993_not
g5266 not n3010 ; n3010_not
g5267 not n3011 ; n3011_not
g5268 not n2988 ; n2988_not
g5269 not n3013 ; n3013_not
g5270 not n3014 ; n3014_not
g5271 not n3008 ; n3008_not
g5272 not n3015 ; n3015_not
g5273 not n3007 ; n3007_not
g5274 not n1883 ; n1883_not
g5275 not n3018 ; n3018_not
g5276 not n3017 ; n3017_not
g5277 not n1890 ; n1890_not
g5278 not n3021 ; n3021_not
g5279 not n1888 ; n1888_not
g5280 not n1861 ; n1861_not
g5281 not n1854 ; n1854_not
g5282 not n3024 ; n3024_not
g5283 not n1832 ; n1832_not
g5284 not n1835 ; n1835_not
g5285 not n1831 ; n1831_not
g5286 not n1850 ; n1850_not
g5287 not n3030 ; n3030_not
g5288 not n3031 ; n3031_not
g5289 not n1845 ; n1845_not
g5290 not n3033 ; n3033_not
g5291 not n3034 ; n3034_not
g5292 not n3028 ; n3028_not
g5293 not n3035 ; n3035_not
g5294 not n3027 ; n3027_not
g5295 not n1818 ; n1818_not
g5296 not n3038 ; n3038_not
g5297 not n3037 ; n3037_not
g5298 not n1825 ; n1825_not
g5299 not n3041 ; n3041_not
g5300 not n1823 ; n1823_not
g5301 not n1796 ; n1796_not
g5302 not n3045 ; n3045_not
g5303 not n3046 ; n3046_not
g5304 not n3048 ; n3048_not
g5305 not n3049 ; n3049_not
g5306 not n3050 ; n3050_not
g5307 not n3052 ; n3052_not
g5308 not n3053 ; n3053_not
g5309 not n3055 ; n3055_not
g5310 not n3056 ; n3056_not
g5311 not n3054 ; n3054_not
g5312 not n3051 ; n3051_not
g5313 not n3058 ; n3058_not
g5314 not n3060 ; n3060_not
g5315 not n3061 ; n3061_not
g5316 not n3063 ; n3063_not
g5317 not n3064 ; n3064_not
g5318 not n3065 ; n3065_not
g5319 not n3067 ; n3067_not
g5320 not n3068 ; n3068_not
g5321 not n3070 ; n3070_not
g5322 not n3071 ; n3071_not
g5323 not n3069 ; n3069_not
g5324 not n3066 ; n3066_not
g5325 not n3073 ; n3073_not
g5326 not n3044 ; n3044_not
g5327 not n3047 ; n3047_not
g5328 not n3072 ; n3072_not
g5329 not n3062 ; n3062_not
g5330 not n3079 ; n3079_not
g5331 not n3080 ; n3080_not
g5332 not n3057 ; n3057_not
g5333 not n3082 ; n3082_not
g5334 not n3083 ; n3083_not
g5335 not n3077 ; n3077_not
g5336 not n3084 ; n3084_not
g5337 not n3076 ; n3076_not
g5338 not n3087 ; n3087_not
g5339 not n3088 ; n3088_not
g5340 not n3090 ; n3090_not
g5341 not n3091 ; n3091_not
g5342 not n3092 ; n3092_not
g5343 not n1213 ; n1213_not
g5344 not n3095 ; n3095_not
g5345 not n3096 ; n3096_not
g5346 not n3098 ; n3098_not
g5347 not n3099 ; n3099_not
g5348 not n3100 ; n3100_not
g5349 not n3102 ; n3102_not
g5350 not n3103 ; n3103_not
g5351 not n3105 ; n3105_not
g5352 not n3106 ; n3106_not
g5353 not n3107 ; n3107_not
g5354 not n3101 ; n3101_not
g5355 not n3108 ; n3108_not
g5356 not n3094 ; n3094_not
g5357 not n3093 ; n3093_not
g5358 not n3086 ; n3086_not
g5359 not n3089 ; n3089_not
g5360 not n3104 ; n3104_not
g5361 not n3113 ; n3113_not
g5362 not n3114 ; n3114_not
g5363 not n3115 ; n3115_not
g5364 not n3097 ; n3097_not
g5365 not n3116 ; n3116_not
g5366 not n3117 ; n3117_not
g5367 not n3118 ; n3118_not
g5368 not n3112 ; n3112_not
g5369 not n3119 ; n3119_not
g5370 not n1785 ; n1785_not
g5371 not n2503 ; n2503_not
g5372 not address[1] ; address[1]_not
g5373 not n3122 ; n3122_not
g5374 not n3123 ; n3123_not
g5375 not n2508 ; n2508_not
g5376 not n3125 ; n3125_not
g5377 not n3126 ; n3126_not
g5378 not n3128 ; n3128_not
g5379 not n3129 ; n3129_not
g5380 not n3131 ; n3131_not
g5381 not n3132 ; n3132_not
g5382 not n2484 ; n2484_not
g5383 not n3134 ; n3134_not
g5384 not n3135 ; n3135_not
g5385 not n2478 ; n2478_not
g5386 not n3137 ; n3137_not
g5387 not n3138 ; n3138_not
g5388 not n2472 ; n2472_not
g5389 not n3140 ; n3140_not
g5390 not n3141 ; n3141_not
g5391 not n3143 ; n3143_not
g5392 not n3144 ; n3144_not
g5393 not n2462 ; n2462_not
g5394 not n3146 ; n3146_not
g5395 not n3147 ; n3147_not
g5396 not n2459 ; n2459_not
g5397 not n3149 ; n3149_not
g5398 not n3150 ; n3150_not
g5399 not n3152 ; n3152_not
g5400 not n3153 ; n3153_not
g5401 not n3155 ; n3155_not
g5402 not n3156 ; n3156_not
g5403 not n3158 ; n3158_not
g5404 not n3159 ; n3159_not
g5405 not n3161 ; n3161_not
g5406 not n3162 ; n3162_not
g5407 not n3164 ; n3164_not
g5408 not n3165 ; n3165_not
g5409 not n3167 ; n3167_not
g5410 not n3168 ; n3168_not
g5411 not n2414 ; n2414_not
g5412 not n3170 ; n3170_not
g5413 not n3171 ; n3171_not
g5414 not n2411 ; n2411_not
g5415 not n3173 ; n3173_not
g5416 not n3174 ; n3174_not
g5417 not n3176 ; n3176_not
g5418 not n3177 ; n3177_not
g5419 not n3179 ; n3179_not
g5420 not n3180 ; n3180_not
g5421 not n3182 ; n3182_not
g5422 not n3183 ; n3183_not
g5423 not n3185 ; n3185_not
g5424 not n3186 ; n3186_not
g5425 not n3188 ; n3188_not
g5426 not n3189 ; n3189_not
g5427 not n3191 ; n3191_not
g5428 not n3192 ; n3192_not
g5429 not n2366 ; n2366_not
g5430 not n3194 ; n3194_not
g5431 not n3195 ; n3195_not
g5432 not n2363 ; n2363_not
g5433 not n3197 ; n3197_not
g5434 not n3198 ; n3198_not
g5435 not n3200 ; n3200_not
g5436 not n3201 ; n3201_not
g5437 not n3203 ; n3203_not
g5438 not n3204 ; n3204_not
g5439 not n3206 ; n3206_not
g5440 not n3207 ; n3207_not
g5441 not n3209 ; n3209_not
g5442 not n3210 ; n3210_not
g5443 not n3212 ; n3212_not
g5444 not n3213 ; n3213_not
g5445 not n3215 ; n3215_not
g5446 not n3216 ; n3216_not
g5447 not n3218 ; n3218_not
g5448 not n3219 ; n3219_not
g5449 not n3221 ; n3221_not
g5450 not n3222 ; n3222_not
g5451 not n3224 ; n3224_not
g5452 not n3225 ; n3225_not
g5453 not n3227 ; n3227_not
g5454 not n3228 ; n3228_not
g5455 not n3230 ; n3230_not
g5456 not n3231 ; n3231_not
g5457 not n3233 ; n3233_not
g5458 not n3234 ; n3234_not
g5459 not n3236 ; n3236_not
g5460 not n3237 ; n3237_not
g5461 not n3239 ; n3239_not
g5462 not n3240 ; n3240_not
g5463 not n3242 ; n3242_not
g5464 not n3243 ; n3243_not
g5465 not n3245 ; n3245_not
g5466 not n3246 ; n3246_not
g5467 not n3248 ; n3248_not
g5468 not n3249 ; n3249_not
g5469 not n3251 ; n3251_not
g5470 not n3252 ; n3252_not
g5471 not n3254 ; n3254_not
g5472 not n3255 ; n3255_not
g5473 not n3257 ; n3257_not
g5474 not n3258 ; n3258_not
g5475 not n3260 ; n3260_not
g5476 not n3261 ; n3261_not
g5477 not n3263 ; n3263_not
g5478 not n3264 ; n3264_not
g5479 not n3266 ; n3266_not
g5480 not n3267 ; n3267_not
g5481 not n3269 ; n3269_not
g5482 not n3270 ; n3270_not
g5483 not n3272 ; n3272_not
g5484 not n3273 ; n3273_not
g5485 not n3275 ; n3275_not
g5486 not n3276 ; n3276_not
g5487 not n3278 ; n3278_not
g5488 not n3279 ; n3279_not
g5489 not n3281 ; n3281_not
g5490 not n3282 ; n3282_not
g5491 not n3284 ; n3284_not
g5492 not n3285 ; n3285_not
g5493 not n3287 ; n3287_not
g5494 not n3288 ; n3288_not
g5495 not n3290 ; n3290_not
g5496 not n3291 ; n3291_not
g5497 not n3293 ; n3293_not
g5498 not n3294 ; n3294_not
g5499 not n3296 ; n3296_not
g5500 not n3297 ; n3297_not
g5501 not n3299 ; n3299_not
g5502 not n3300 ; n3300_not
g5503 not n3302 ; n3302_not
g5504 not n3303 ; n3303_not
g5505 not n3305 ; n3305_not
g5506 not n3306 ; n3306_not
g5507 not n3308 ; n3308_not
g5508 not n3309 ; n3309_not
g5509 not n3311 ; n3311_not
g5510 not n3312 ; n3312_not
g5511 not n3314 ; n3314_not
g5512 not n3315 ; n3315_not
g5513 not n3317 ; n3317_not
g5514 not n3318 ; n3318_not
g5515 not n3320 ; n3320_not
g5516 not n3321 ; n3321_not
g5517 not n3323 ; n3323_not
g5518 not n3324 ; n3324_not
g5519 not n3326 ; n3326_not
g5520 not n3327 ; n3327_not
g5521 not n3329 ; n3329_not
g5522 not n3330 ; n3330_not
g5523 not n3332 ; n3332_not
g5524 not n3333 ; n3333_not
g5525 not n3335 ; n3335_not
g5526 not n3336 ; n3336_not
g5527 not n3338 ; n3338_not
g5528 not n3339 ; n3339_not
g5529 not n3341 ; n3341_not
g5530 not n3342 ; n3342_not
g5531 not n3344 ; n3344_not
g5532 not n3345 ; n3345_not
g5533 not n3347 ; n3347_not
g5534 not n3348 ; n3348_not
g5535 not n3350 ; n3350_not
g5536 not n3351 ; n3351_not
g5537 not n3353 ; n3353_not
g5538 not n3354 ; n3354_not
g5539 not n3356 ; n3356_not
g5540 not n3357 ; n3357_not
g5541 not n3359 ; n3359_not
g5542 not n3360 ; n3360_not
g5543 not n3362 ; n3362_not
g5544 not n3363 ; n3363_not
g5545 not n3365 ; n3365_not
g5546 not n3366 ; n3366_not
g5547 not n3368 ; n3368_not
g5548 not n3369 ; n3369_not
g5549 not n3371 ; n3371_not
g5550 not n3372 ; n3372_not
g5551 not n3374 ; n3374_not
g5552 not n3375 ; n3375_not
g5553 not n3377 ; n3377_not
g5554 not n3378 ; n3378_not
g5555 not n3380 ; n3380_not
g5556 not n3381 ; n3381_not
g5557 not n3383 ; n3383_not
g5558 not n3384 ; n3384_not
g5559 not n3386 ; n3386_not
g5560 not n3387 ; n3387_not
g5561 not n3389 ; n3389_not
g5562 not n3390 ; n3390_not
g5563 not n3392 ; n3392_not
g5564 not n3393 ; n3393_not
g5565 not n3395 ; n3395_not
g5566 not n3396 ; n3396_not
g5567 not n3398 ; n3398_not
g5568 not n3399 ; n3399_not
g5569 not n3401 ; n3401_not
g5570 not n3402 ; n3402_not
g5571 not n3404 ; n3404_not
g5572 not n3405 ; n3405_not
g5573 not n3407 ; n3407_not
g5574 not n3408 ; n3408_not
g5575 not n3410 ; n3410_not
g5576 not n3411 ; n3411_not
g5577 not n3413 ; n3413_not
g5578 not n3414 ; n3414_not
g5579 not n3416 ; n3416_not
g5580 not n3417 ; n3417_not
g5581 not n3419 ; n3419_not
g5582 not n3420 ; n3420_not
g5583 not n3422 ; n3422_not
g5584 not n3423 ; n3423_not
g5585 not n3425 ; n3425_not
g5586 not n3426 ; n3426_not
g5587 not n3428 ; n3428_not
g5588 not n3429 ; n3429_not
g5589 not n3431 ; n3431_not
g5590 not n3432 ; n3432_not
g5591 not n3434 ; n3434_not
g5592 not n3435 ; n3435_not
g5593 not n3437 ; n3437_not
g5594 not n3438 ; n3438_not
g5595 not n3440 ; n3440_not
g5596 not n3441 ; n3441_not
g5597 not n3443 ; n3443_not
g5598 not n3444 ; n3444_not
g5599 not n3446 ; n3446_not
g5600 not n3447 ; n3447_not
g5601 not n3449 ; n3449_not
g5602 not n3450 ; n3450_not
g5603 not n3452 ; n3452_not
g5604 not n3453 ; n3453_not
g5605 not n3455 ; n3455_not
g5606 not n3456 ; n3456_not
g5607 not n3458 ; n3458_not
g5608 not n3459 ; n3459_not
g5609 not n3461 ; n3461_not
g5610 not n3462 ; n3462_not
g5611 not n3464 ; n3464_not
g5612 not n3465 ; n3465_not
g5613 not n3467 ; n3467_not
g5614 not n3468 ; n3468_not
g5615 not n3470 ; n3470_not
g5616 not n3471 ; n3471_not
g5617 not n3473 ; n3473_not
g5618 not n3474 ; n3474_not
g5619 not n3476 ; n3476_not
g5620 not n3477 ; n3477_not
g5621 not n3479 ; n3479_not
g5622 not n3480 ; n3480_not
g5623 not n3482 ; n3482_not
g5624 not n3483 ; n3483_not
g5625 not n3485 ; n3485_not
g5626 not n3486 ; n3486_not
g5627 not n3488 ; n3488_not
g5628 not n3489 ; n3489_not
g5629 not n3491 ; n3491_not
g5630 not n3492 ; n3492_not
g5631 not n3494 ; n3494_not
g5632 not n3495 ; n3495_not
g5633 not n3497 ; n3497_not
g5634 not n3498 ; n3498_not
g5635 not n3500 ; n3500_not
g5636 not n3501 ; n3501_not
g5637 not n3503 ; n3503_not
g5638 not n3505 ; n3505_not
g5639 not n3506 ; n3506_not
o result[0]
o result[1]
o result[2]
o result[3]
o result[4]
o result[5]
o result[6]
o result[7]
o result[8]
o result[9]
o result[10]
o result[11]
o result[12]
o result[13]
o result[14]
o result[15]
o result[16]
o result[17]
o result[18]
o result[19]
o result[20]
o result[21]
o result[22]
o result[23]
o result[24]
o result[25]
o result[26]
o result[27]
o result[28]
o result[29]
o result[30]
o result[31]
o result[32]
o result[33]
o result[34]
o result[35]
o result[36]
o result[37]
o result[38]
o result[39]
o result[40]
o result[41]
o result[42]
o result[43]
o result[44]
o result[45]
o result[46]
o result[47]
o result[48]
o result[49]
o result[50]
o result[51]
o result[52]
o result[53]
o result[54]
o result[55]
o result[56]
o result[57]
o result[58]
o result[59]
o result[60]
o result[61]
o result[62]
o result[63]
o result[64]
o result[65]
o result[66]
o result[67]
o result[68]
o result[69]
o result[70]
o result[71]
o result[72]
o result[73]
o result[74]
o result[75]
o result[76]
o result[77]
o result[78]
o result[79]
o result[80]
o result[81]
o result[82]
o result[83]
o result[84]
o result[85]
o result[86]
o result[87]
o result[88]
o result[89]
o result[90]
o result[91]
o result[92]
o result[93]
o result[94]
o result[95]
o result[96]
o result[97]
o result[98]
o result[99]
o result[100]
o result[101]
o result[102]
o result[103]
o result[104]
o result[105]
o result[106]
o result[107]
o result[108]
o result[109]
o result[110]
o result[111]
o result[112]
o result[113]
o result[114]
o result[115]
o result[116]
o result[117]
o result[118]
o result[119]
o result[120]
o result[121]
o result[122]
o result[123]
o result[124]
o result[125]
o result[126]
o result[127]
o address[0]
