name sin
i a[0]
i a[1]
i a[2]
i a[3]
i a[4]
i a[5]
i a[6]
i a[7]
i a[8]
i a[9]
i a[10]
i a[11]
i a[12]
i a[13]
i a[14]
i a[15]
i a[16]
i a[17]
i a[18]
i a[19]
i a[20]
i a[21]
i a[22]
i a[23]

o sin[0]
o sin[1]
o sin[2]
o sin[3]
o sin[4]
o sin[5]
o sin[6]
o sin[7]
o sin[8]
o sin[9]
o sin[10]
o sin[11]
o sin[12]
o sin[13]
o sin[14]
o sin[15]
o sin[16]
o sin[17]
o sin[18]
o sin[19]
o sin[20]
o sin[21]
o sin[22]
o sin[23]
o sin[24]

g1 and a[21] a[22] ; n50
g2 nor a[1] a[2] ; n51
g3 and a[0]_not n51 ; n52
g4 and a[3]_not n52 ; n53
g5 and a[4]_not n53 ; n54
g6 and a[5]_not n54 ; n55
g7 and a[6]_not n55 ; n56
g8 and a[7]_not n56 ; n57
g9 and a[8]_not n57 ; n58
g10 and a[9]_not n58 ; n59
g11 and a[10]_not n59 ; n60
g12 and a[11]_not n60 ; n61
g13 and a[12]_not n61 ; n62
g14 and a[13]_not n62 ; n63
g15 and a[14]_not n63 ; n64
g16 and a[15]_not n64 ; n65
g17 and a[16]_not n65 ; n66
g18 and a[17]_not n66 ; n67
g19 and a[18]_not n67 ; n68
g20 and a[19]_not n68 ; n69
g21 and a[20]_not n69 ; n70
g22 and a[21]_not n70 ; n71
g23 and a[21] n70_not ; n72
g24 nor n71 n72 ; n73
g25 and a[22]_not n73 ; n74
g26 nor n50 n74 ; n75
g27 and a[20] a[22] ; n76
g28 and a[20] n69_not ; n77
g29 nor n70 n77 ; n78
g30 and a[22]_not n78 ; n79
g31 nor n76 n79 ; n80
g32 and n75 n80 ; n81
g33 and a[15] a[22] ; n82
g34 nor a[22] n65 ; n83
g35 and a[15] n64_not ; n84
g36 and n83 n84_not ; n85
g37 nor n82 n85 ; n86
g38 and n81 n86 ; n87
g39 nor a[22] n68 ; n88
g40 and a[19] n88_not ; n89
g41 and a[19]_not n88 ; n90
g42 nor n89 n90 ; n91
g43 and a[18] a[22] ; n92
g44 and a[18] n67_not ; n93
g45 and n88 n93_not ; n94
g46 nor n92 n94 ; n95
g47 nor n91 n95 ; n96
g48 nor a[22] n66 ; n97
g49 and a[17] n97_not ; n98
g50 and a[17]_not n97 ; n99
g51 nor n98 n99 ; n100
g52 and a[16] n83_not ; n101
g53 and a[16]_not n83 ; n102
g54 nor n101 n102 ; n103
g55 and n100_not n103 ; n104
g56 and n96 n104 ; n105
g57 and n87 n105 ; n106
g58 and n100 n103 ; n107
g59 and n96 n107 ; n108
g60 and n75 n80_not ; n109
g61 and n86 n109 ; n110
g62 and n108 n110 ; n111
g63 and n91_not n95 ; n112
g64 and n107 n112 ; n113
g65 and n110 n113 ; n114
g66 and n86_not n109 ; n115
g67 and n91 n95_not ; n116
g68 and n107 n116 ; n117
g69 and n115 n117 ; n118
g70 and n75_not n80 ; n119
g71 and n86_not n119 ; n120
g72 and n100 n103_not ; n121
g73 and n112 n121 ; n122
g74 and n120 n122 ; n123
g75 nor n75 n80 ; n124
g76 and n86_not n124 ; n125
g77 and n104 n112 ; n126
g78 and n125 n126 ; n127
g79 and n86 n124 ; n128
g80 and n105 n128 ; n129
g81 and n81 n86_not ; n130
g82 and n104 n116 ; n131
g83 and n130 n131 ; n132
g84 and n105 n120 ; n133
g85 and n122 n125 ; n134
g86 nor n100 n103 ; n135
g87 and n116 n135 ; n136
g88 and n125 n136 ; n137
g89 and n128 n136 ; n138
g90 and n122 n128 ; n139
g91 and n128 n131 ; n140
g92 nor n139 n140 ; n141
g93 and n105 n110 ; n142
g94 and n96 n121 ; n143
g95 and n128 n143 ; n144
g96 nor n142 n144 ; n145
g97 and n105 n115 ; n146
g98 and n116 n121 ; n147
g99 and n110 n147 ; n148
g100 nor n146 n148 ; n149
g101 and n126 n128 ; n150
g102 and n112 n135 ; n151
g103 and n128 n151 ; n152
g104 nor n150 n152 ; n153
g105 and n130 n136 ; n154
g106 and n105 n125 ; n155
g107 nor n154 n155 ; n156
g108 and n153 n156 ; n157
g109 and n149 n157 ; n158
g110 and n145 n158 ; n159
g111 and n141 n159 ; n160
g112 and n138_not n160 ; n161
g113 and n137_not n161 ; n162
g114 and n134_not n162 ; n163
g115 and n133_not n163 ; n164
g116 and n132_not n164 ; n165
g117 and n110 n143 ; n166
g118 and n120 n151 ; n167
g119 and n87 n151 ; n168
g120 and n115 n122 ; n169
g121 and n91 n95 ; n170
g122 and n107 n170 ; n171
g123 and n115 n171 ; n172
g124 and n86 n119 ; n173
g125 and n151 n173 ; n174
g126 and n108 n125 ; n175
g127 and n125 n143 ; n176
g128 and n117 n173 ; n177
g129 and n108 n128 ; n178
g130 nor n177 n178 ; n179
g131 and n176_not n179 ; n180
g132 and n175_not n180 ; n181
g133 and n174_not n181 ; n182
g134 and n172_not n182 ; n183
g135 and n169_not n183 ; n184
g136 and n168_not n184 ; n185
g137 and n108 n120 ; n186
g138 and n135 n170 ; n187
g139 and n128 n187 ; n188
g140 nor n186 n188 ; n189
g141 and n110 n151 ; n190
g142 and n117 n120 ; n191
g143 and n120 n126 ; n192
g144 and n121 n170 ; n193
g145 and n125 n193 ; n194
g146 and n96 n135 ; n195
g147 and n128 n195 ; n196
g148 nor n194 n196 ; n197
g149 and n192_not n197 ; n198
g150 and n191_not n198 ; n199
g151 and n190_not n199 ; n200
g152 and n189 n200 ; n201
g153 and n185 n201 ; n202
g154 and n167_not n202 ; n203
g155 and n166_not n203 ; n204
g156 and n104 n170 ; n205
g157 and n115 n205 ; n206
g158 and n120 n131 ; n207
g159 and n128 n147 ; n208
g160 nor n207 n208 ; n209
g161 and n206_not n209 ; n210
g162 and n130 n147 ; n211
g163 and n115 n195 ; n212
g164 and n171 n173 ; n213
g165 and n125 n171 ; n214
g166 and n117 n130 ; n215
g167 and n110 n126 ; n216
g168 and n120 n147 ; n217
g169 and n108 n173 ; n218
g170 and n125 n187 ; n219
g171 and n125 n131 ; n220
g172 and n125 n147 ; n221
g173 and n128 n193 ; n222
g174 and n122 n130 ; n223
g175 and n115 n126 ; n224
g176 and n120 n143 ; n225
g177 and n105 n173 ; n226
g178 and n125 n151 ; n227
g179 and n113 n125 ; n228
g180 nor n227 n228 ; n229
g181 and n226_not n229 ; n230
g182 and n225_not n230 ; n231
g183 and n224_not n231 ; n232
g184 and n223_not n232 ; n233
g185 and n115 n187 ; n234
g186 and n105 n130 ; n235
g187 nor n234 n235 ; n236
g188 and n130 n187 ; n237
g189 and n130 n205 ; n238
g190 nor n237 n238 ; n239
g191 and n236 n239 ; n240
g192 and n233 n240 ; n241
g193 and n222_not n241 ; n242
g194 and n221_not n242 ; n243
g195 and n220_not n243 ; n244
g196 and n219_not n244 ; n245
g197 and n218_not n245 ; n246
g198 and n217_not n246 ; n247
g199 and n216_not n247 ; n248
g200 and n215_not n248 ; n249
g201 and n214_not n249 ; n250
g202 and n213_not n250 ; n251
g203 and n212_not n251 ; n252
g204 and n211_not n252 ; n253
g205 and n173 n193 ; n254
g206 and n120 n195 ; n255
g207 nor n254 n255 ; n256
g208 and n113 n173 ; n257
g209 and n87 n193 ; n258
g210 nor n257 n258 ; n259
g211 and n256 n259 ; n260
g212 and n253 n260 ; n261
g213 and n210 n261 ; n262
g214 and n204 n262 ; n263
g215 and n165 n263 ; n264
g216 and n129_not n264 ; n265
g217 and n127_not n265 ; n266
g218 and n123_not n266 ; n267
g219 and n118_not n267 ; n268
g220 and n114_not n268 ; n269
g221 and n111_not n269 ; n270
g222 and n106_not n270 ; n271
g223 nor a[22] n54 ; n272
g224 and a[5] n272_not ; n273
g225 and a[5]_not n272 ; n274
g226 nor n273 n274 ; n275
g227 and a[4] a[22] ; n276
g228 and a[4] n53_not ; n277
g229 and n272 n277_not ; n278
g230 nor n276 n278 ; n279
g231 and n275 n279_not ; n280
g232 and n275_not n279 ; n281
g233 nor n280 n281 ; n282
g234 nor a[22] n52 ; n283
g235 and a[3] n283_not ; n284
g236 and a[3]_not n283 ; n285
g237 nor n284 n285 ; n286
g238 and a[2] a[22] ; n287
g239 nor a[0] a[1] ; n288
g240 and a[2] n288_not ; n289
g241 and n283 n289_not ; n290
g242 nor n287 n290 ; n291
g243 and n286 n291_not ; n292
g244 and n286_not n291 ; n293
g245 nor n292 n293 ; n294
g246 and n282 n294_not ; n295
g247 and n130 n151 ; n296
g248 and n108 n115 ; n297
g249 and n113 n115 ; n298
g250 and n122 n173 ; n299
g251 and n120 n205 ; n300
g252 nor n211 n300 ; n301
g253 and n115 n131 ; n302
g254 nor n111 n302 ; n303
g255 and n179 n303 ; n304
g256 and n301 n304 ; n305
g257 and n137_not n305 ; n306
g258 and n299_not n306 ; n307
g259 and n191_not n307 ; n308
g260 and n298_not n308 ; n309
g261 and n297_not n309 ; n310
g262 and n296_not n310 ; n311
g263 and n173 n195 ; n312
g264 and n120 n136 ; n313
g265 nor n221 n313 ; n314
g266 and n110 n187 ; n315
g267 nor n114 n315 ; n316
g268 and n125 n205 ; n317
g269 nor n129 n317 ; n318
g270 and n207_not n318 ; n319
g271 and n316 n319 ; n320
g272 and n314 n320 ; n321
g273 and n312_not n321 ; n322
g274 and n212_not n322 ; n323
g275 and n87 n171 ; n324
g276 nor n123 n324 ; n325
g277 and n87 n147 ; n326
g278 and n136 n173 ; n327
g279 and n128 n205 ; n328
g280 and n147 n173 ; n329
g281 nor n328 n329 ; n330
g282 and n255_not n330 ; n331
g283 and n327_not n331 ; n332
g284 and n168_not n332 ; n333
g285 and n326_not n333 ; n334
g286 and n110 n193 ; n335
g287 and n113 n120 ; n336
g288 and n113 n128 ; n337
g289 nor n188 n337 ; n338
g290 and n175_not n338 ; n339
g291 and n336_not n339 ; n340
g292 and n335_not n340 ; n341
g293 and n108 n130 ; n342
g294 and n173 n187 ; n343
g295 nor n342 n343 ; n344
g296 and n130 n171 ; n345
g297 nor n150 n345 ; n346
g298 and n110 n195 ; n347
g299 and n131 n173 ; n348
g300 nor n347 n348 ; n349
g301 and n126 n173 ; n350
g302 and n87 n113 ; n351
g303 nor n192 n226 ; n352
g304 and n351_not n352 ; n353
g305 and n217_not n353 ; n354
g306 and n216_not n354 ; n355
g307 and n110 n171 ; n356
g308 and n110 n136 ; n357
g309 and n110 n205 ; n358
g310 and n110 n117 ; n359
g311 and n120 n187 ; n360
g312 and n115 n147 ; n361
g313 nor n360 n361 ; n362
g314 and n359_not n362 ; n363
g315 and n358_not n363 ; n364
g316 and n357_not n364 ; n365
g317 and n356_not n365 ; n366
g318 and n87 n195 ; n367
g319 and n87 n126 ; n368
g320 nor n127 n368 ; n369
g321 and n173 n205 ; n370
g322 and n369 n370_not ; n371
g323 and n367_not n371 ; n372
g324 nor n106 n215 ; n373
g325 and n372 n373 ; n374
g326 and n366 n374 ; n375
g327 and n355 n375 ; n376
g328 and n174_not n376 ; n377
g329 and n133_not n377 ; n378
g330 and n146_not n378 ; n379
g331 and n223_not n379 ; n380
g332 and n156 n380 ; n381
g333 and n350_not n381 ; n382
g334 and n349 n382 ; n383
g335 and n346 n383 ; n384
g336 and n259 n384 ; n385
g337 and n344 n385 ; n386
g338 and n341 n386 ; n387
g339 and n334 n387 ; n388
g340 and n325 n388 ; n389
g341 and n323 n389 ; n390
g342 and n311 n390 ; n391
g343 and n208_not n391 ; n392
g344 and n134_not n392 ; n393
g345 and n125 n195 ; n394
g346 nor n192 n350 ; n395
g347 nor n174 n337 ; n396
g348 nor n207 n327 ; n397
g349 and n396 n397 ; n398
g350 and n314 n398 ; n399
g351 and n141 n399 ; n400
g352 and n208_not n400 ; n401
g353 and n228_not n401 ; n402
g354 and n395 n402 ; n403
g355 and n167_not n403 ; n404
g356 and n117 n125 ; n405
g357 nor n137 n257 ; n406
g358 and n336_not n406 ; n407
g359 and n117 n128 ; n408
g360 nor n138 n408 ; n409
g361 and n220_not n409 ; n410
g362 and n299_not n410 ; n411
g363 and n407 n411 ; n412
g364 and n405_not n412 ; n413
g365 and n123_not n413 ; n414
g366 and n128 n171 ; n415
g367 nor n255 n415 ; n416
g368 and n143 n173 ; n417
g369 and n153 n189 ; n418
g370 and n127_not n418 ; n419
g371 and n219_not n419 ; n420
g372 and n225_not n420 ; n421
g373 and n417_not n421 ; n422
g374 and n218_not n422 ; n423
g375 and n416 n423 ; n424
g376 and n414 n424 ; n425
g377 and n222_not n425 ; n426
g378 and n144_not n426 ; n427
g379 and n129_not n427 ; n428
g380 and n176_not n428 ; n429
g381 and n214_not n429 ; n430
g382 and n134_not n430 ; n431
g383 nor n155 n194 ; n432
g384 nor n178 n227 ; n433
g385 and n175_not n433 ; n434
g386 and n312_not n434 ; n435
g387 and n226_not n435 ; n436
g388 and n133_not n436 ; n437
g389 and n432 n437 ; n438
g390 and n431 n438 ; n439
g391 and n404 n439 ; n440
g392 and n328_not n440 ; n441
g393 and n196_not n441 ; n442
g394 and n317_not n442 ; n443
g395 and n394_not n443 ; n444
g396 and n87 n122 ; n445
g397 and n120 n171 ; n446
g398 and n115 n151 ; n447
g399 nor n190 n447 ; n448
g400 and n115 n143 ; n449
g401 nor n297 n449 ; n450
g402 and n166_not n450 ; n451
g403 and n448 n451 ; n452
g404 and n146_not n452 ; n453
g405 nor n254 n343 ; n454
g406 and n224_not n454 ; n455
g407 and n212_not n455 ; n456
g408 and n142_not n456 ; n457
g409 and n120 n193 ; n458
g410 nor n300 n458 ; n459
g411 nor n360 n370 ; n460
g412 and n349 n460 ; n461
g413 and n459 n461 ; n462
g414 and n457 n462 ; n463
g415 and n453 n463 ; n464
g416 and n213_not n464 ; n465
g417 and n446_not n465 ; n466
g418 and n111_not n466 ; n467
g419 and n113 n130 ; n468
g420 and n126 n130 ; n469
g421 and n87 n108 ; n470
g422 and n130 n195 ; n471
g423 and n87 n143 ; n472
g424 nor n177 n329 ; n473
g425 nor n235 n356 ; n474
g426 nor n191 n217 ; n475
g427 and n172_not n475 ; n476
g428 and n130 n143 ; n477
g429 nor n342 n477 ; n478
g430 and n476 n478 ; n479
g431 and n474 n479 ; n480
g432 and n473 n480 ; n481
g433 and n106_not n481 ; n482
g434 and n367_not n482 ; n483
g435 and n472_not n483 ; n484
g436 and n471_not n484 ; n485
g437 and n470_not n485 ; n486
g438 and n168_not n486 ; n487
g439 and n296_not n487 ; n488
g440 and n469_not n488 ; n489
g441 and n468_not n489 ; n490
g442 and n467 n490 ; n491
g443 and n368_not n491 ; n492
g444 and n445_not n492 ; n493
g445 and n223_not n493 ; n494
g446 and n115 n193 ; n495
g447 nor n118 n335 ; n496
g448 and n495_not n496 ; n497
g449 and n358_not n497 ; n498
g450 and n315_not n498 ; n499
g451 and n234_not n499 ; n500
g452 and n206_not n500 ; n501
g453 and n359_not n501 ; n502
g454 and n110 n122 ; n503
g455 and n115 n136 ; n504
g456 nor n216 n504 ; n505
g457 and n110 n131 ; n506
g458 nor n357 n361 ; n507
g459 and n506_not n507 ; n508
g460 and n505 n508 ; n509
g461 and n302_not n509 ; n510
g462 and n298_not n510 ; n511
g463 and n169_not n511 ; n512
g464 and n114_not n512 ; n513
g465 and n503_not n513 ; n514
g466 and n467 n514 ; n515
g467 and n475 n515 ; n516
g468 and n473 n516 ; n517
g469 and n502 n517 ; n518
g470 and n148_not n518 ; n519
g471 nor n494 n519 ; n520
g472 and a[14] a[22] ; n521
g473 and a[14] n63_not ; n522
g474 nor n64 n522 ; n523
g475 and a[22]_not n523 ; n524
g476 nor n521 n524 ; n525
g477 nor a[22] n62 ; n526
g478 and a[13] n526_not ; n527
g479 and a[13]_not n526 ; n528
g480 nor n527 n528 ; n529
g481 and n525_not n529 ; n530
g482 and n525 n529_not ; n531
g483 nor n530 n531 ; n532
g484 and n520 n532 ; n533
g485 nor n520 n532 ; n534
g486 nor n533 n534 ; n535
g487 and n444_not n535 ; n536
g488 and n494 n519_not ; n537
g489 and n494_not n519 ; n538
g490 nor n537 n538 ; n539
g491 and n494 n519 ; n540
g492 and n444 n540_not ; n541
g493 and n539 n541_not ; n542
g494 and n525_not n542 ; n543
g495 nor n444 n520 ; n544
g496 nor n539 n544 ; n545
g497 and n525 n544_not ; n546
g498 nor n545 n546 ; n547
g499 and n543_not n547 ; n548
g500 nor n444 n529 ; n549
g501 and n548 n549_not ; n550
g502 and n548_not n549 ; n551
g503 and n87 n136 ; n552
g504 and n87 n205 ; n553
g505 and n87 n131 ; n554
g506 nor n238 n554 ; n555
g507 and n208_not n555 ; n556
g508 and n221_not n556 ; n557
g509 and n367_not n557 ; n558
g510 nor n225 n417 ; n559
g511 and n296_not n559 ; n560
g512 nor n234 n471 ; n561
g513 and n237_not n561 ; n562
g514 nor n227 n394 ; n563
g515 and n127_not n563 ; n564
g516 and n562 n564 ; n565
g517 and n560 n565 ; n566
g518 and n558 n566 ; n567
g519 and n185 n567 ; n568
g520 and n129_not n568 ; n569
g521 and n348_not n569 ; n570
g522 and n553_not n570 ; n571
g523 nor n167 n220 ; n572
g524 and n191_not n572 ; n573
g525 and n337_not n573 ; n574
g526 and n360_not n574 ; n575
g527 and n212_not n575 ; n576
g528 and n470_not n576 ; n577
g529 nor n118 n196 ; n578
g530 and n114_not n578 ; n579
g531 and n503_not n579 ; n580
g532 and n469_not n580 ; n581
g533 nor n218 n343 ; n582
g534 and n329_not n582 ; n583
g535 and n449_not n583 ; n584
g536 nor n298 n347 ; n585
g537 and n356_not n585 ; n586
g538 and n165 n228_not ; n587
g539 and n359_not n587 ; n588
g540 and n87 n187 ; n589
g541 nor n186 n589 ; n590
g542 and n588 n590 ; n591
g543 and n586 n591 ; n592
g544 and n584 n592 ; n593
g545 and n581 n593 ; n594
g546 and n577 n594 ; n595
g547 and n571 n595 ; n596
g548 and n355 n596 ; n597
g549 and n552_not n597 ; n598
g550 and n87 n117 ; n599
g551 and n141 n373 ; n600
g552 and n220_not n600 ; n601
g553 and n134_not n601 ; n602
g554 and n172_not n602 ; n603
g555 and n298_not n603 ; n604
g556 and n506_not n604 ; n605
g557 and n554_not n605 ; n606
g558 nor n222 n337 ; n607
g559 and n114_not n607 ; n608
g560 nor n317 n405 ; n609
g561 and n474 n609 ; n610
g562 and n227_not n610 ; n611
g563 and n348_not n611 ; n612
g564 and n329_not n612 ; n613
g565 and n154_not n613 ; n614
g566 and n153 n432 ; n615
g567 and n505 n615 ; n616
g568 and n614 n616 ; n617
g569 and n408_not n617 ; n618
g570 and n188_not n618 ; n619
g571 and n129_not n619 ; n620
g572 and n217_not n620 ; n621
g573 and n357_not n621 ; n622
g574 and n326_not n622 ; n623
g575 and n394_not n623 ; n624
g576 and n351_not n624 ; n625
g577 nor n208 n214 ; n626
g578 and n137_not n626 ; n627
g579 and n169_not n627 ; n628
g580 and n625 n628 ; n629
g581 and n344 n629 ; n630
g582 and n608 n630 ; n631
g583 and n606 n631 ; n632
g584 and n191_not n632 ; n633
g585 and n446_not n633 ; n634
g586 and n599_not n634 ; n635
g587 and n211_not n635 ; n636
g588 nor n312 n415 ; n637
g589 nor n176 n503 ; n638
g590 and n637 n638 ; n639
g591 and n196_not n639 ; n640
g592 and n175_not n640 ; n641
g593 and n300_not n641 ; n642
g594 and n302_not n642 ; n643
g595 nor n213 n472 ; n644
g596 nor n138 n228 ; n645
g597 and n477_not n645 ; n646
g598 nor n127 n328 ; n647
g599 and n370_not n647 ; n648
g600 and n256 n648 ; n649
g601 and n144_not n649 ; n650
g602 and n221_not n650 ; n651
g603 and n471_not n651 ; n652
g604 and n132_not n652 ; n653
g605 and n219_not n653 ; n654
g606 and n458_not n654 ; n655
g607 and n179 n655 ; n656
g608 and n646 n656 ; n657
g609 and n644 n657 ; n658
g610 and n643 n658 ; n659
g611 and n636 n659 ; n660
g612 and n362 n660 ; n661
g613 and n552_not n661 ; n662
g614 and n367_not n662 ; n663
g615 nor n598 n663 ; n664
g616 nor n494 n664 ; n665
g617 nor a[22] n60 ; n666
g618 and a[11] n666_not ; n667
g619 and a[11]_not n666 ; n668
g620 nor n667 n668 ; n669
g621 nor n444 n669 ; n670
g622 and n665_not n670 ; n671
g623 and n665 n670_not ; n672
g624 nor n671 n672 ; n673
g625 and a[12] a[22] ; n674
g626 and a[12] n61_not ; n675
g627 and n526 n675_not ; n676
g628 nor n674 n676 ; n677
g629 nor n444 n677 ; n678
g630 and n673 n678 ; n679
g631 nor n671 n679 ; n680
g632 nor n550 n680 ; n681
g633 and n551_not n681 ; n682
g634 nor n550 n682 ; n683
g635 nor n539 n541 ; n684
g636 and n525_not n684 ; n685
g637 and n525 n545 ; n686
g638 and n539 n544_not ; n687
g639 and n529 n687 ; n688
g640 and n529_not n542 ; n689
g641 nor n688 n689 ; n690
g642 and n686_not n690 ; n691
g643 and n685_not n691 ; n692
g644 and n598 n663_not ; n693
g645 and n598_not n663 ; n694
g646 nor n693 n694 ; n695
g647 and n598 n663 ; n696
g648 and n494 n696_not ; n697
g649 and n695 n697_not ; n698
g650 and n525_not n698 ; n699
g651 nor n665 n695 ; n700
g652 and n525 n665_not ; n701
g653 nor n700 n701 ; n702
g654 and n699_not n702 ; n703
g655 and n670_not n703 ; n704
g656 and n529_not n684 ; n705
g657 and n529 n545 ; n706
g658 and n677 n687 ; n707
g659 and n542 n677_not ; n708
g660 nor n707 n708 ; n709
g661 and n706_not n709 ; n710
g662 and n705_not n710 ; n711
g663 and n670 n703_not ; n712
g664 nor n704 n712 ; n713
g665 and n711 n713 ; n714
g666 nor n704 n714 ; n715
g667 and n692 n715_not ; n716
g668 and n692_not n715 ; n717
g669 nor n716 n717 ; n718
g670 nor n673 n678 ; n719
g671 nor n679 n719 ; n720
g672 and n718 n720 ; n721
g673 nor n716 n721 ; n722
g674 nor n680 n682 ; n723
g675 and n551_not n683 ; n724
g676 nor n723 n724 ; n725
g677 and n722_not n725 ; n726
g678 and n722 n725_not ; n727
g679 nor n726 n727 ; n728
g680 nor n222 n415 ; n729
g681 and n219_not n729 ; n730
g682 and n359_not n730 ; n731
g683 and n166_not n731 ; n732
g684 and n470_not n732 ; n733
g685 and n368_not n733 ; n734
g686 and n345_not n734 ; n735
g687 and n130 n193 ; n736
g688 nor n123 n167 ; n737
g689 and n216_not n737 ; n738
g690 and n736_not n738 ; n739
g691 nor n337 n495 ; n740
g692 and n503_not n740 ; n741
g693 and n506_not n741 ; n742
g694 and n351_not n742 ; n743
g695 and n235_not n743 ; n744
g696 and n476 n744 ; n745
g697 and n739 n745 ; n746
g698 and n139_not n746 ; n747
g699 and n504_not n747 ; n748
g700 and n297_not n748 ; n749
g701 and n206_not n749 ; n750
g702 and n106_not n750 ; n751
g703 and n238_not n751 ; n752
g704 nor n132 n298 ; n753
g705 and n348_not n645 ; n754
g706 and n350_not n754 ; n755
g707 and n218_not n755 ; n756
g708 and n148_not n756 ; n757
g709 nor n177 n211 ; n758
g710 and n215_not n758 ; n759
g711 nor n212 n472 ; n760
g712 and n759 n760 ; n761
g713 and n757 n761 ; n762
g714 and n753 n762 ; n763
g715 and n188_not n763 ; n764
g716 and n257_not n764 ; n765
g717 and n142_not n765 ; n766
g718 and n552_not n766 ; n767
g719 and n445_not n767 ; n768
g720 nor n137 n313 ; n769
g721 and n447_not n769 ; n770
g722 and n315_not n770 ; n771
g723 and n168_not n771 ; n772
g724 and n471_not n772 ; n773
g725 nor n214 n405 ; n774
g726 and n302_not n774 ; n775
g727 nor n254 n300 ; n776
g728 and n225_not n776 ; n777
g729 and n775 n777 ; n778
g730 and n773 n778 ; n779
g731 and n768 n779 ; n780
g732 and n752 n780 ; n781
g733 and n735 n781 ; n782
g734 and n408_not n782 ; n783
g735 and n226_not n783 ; n784
g736 and n133_not n784 ; n785
g737 and n237_not n785 ; n786
g738 nor n166 n226 ; n787
g739 and n237_not n787 ; n788
g740 and n477_not n788 ; n789
g741 nor n169 n186 ; n790
g742 and n347_not n790 ; n791
g743 and n223_not n791 ; n792
g744 nor n111 n176 ; n793
g745 and n470_not n793 ; n794
g746 nor n134 n178 ; n795
g747 and n212_not n795 ; n796
g748 and n794 n796 ; n797
g749 and n648 n797 ; n798
g750 and n792 n798 ; n799
g751 and n219_not n799 ; n800
g752 and n350_not n800 ; n801
g753 and n417_not n801 ; n802
g754 and n133_not n802 ; n803
g755 and n315_not n803 ; n804
g756 and n106_not n804 ; n805
g757 nor n225 n299 ; n806
g758 nor n123 n175 ; n807
g759 nor n144 n336 ; n808
g760 nor n458 n589 ; n809
g761 and n301 n809 ; n810
g762 and n149 n810 ; n811
g763 and n258_not n811 ; n812
g764 and n368_not n812 ; n813
g765 and n297_not n813 ; n814
g766 and n206_not n814 ; n815
g767 and n625 n815 ; n816
g768 and n808 n816 ; n817
g769 and n807 n817 ; n818
g770 and n806 n818 ; n819
g771 and n805 n819 ; n820
g772 and n789 n820 ; n821
g773 and n172_not n821 ; n822
g774 and n578 n822 ; n823
g775 and n358_not n823 ; n824
g776 and n736_not n824 ; n825
g777 and n296_not n825 ; n826
g778 nor n786 n826 ; n827
g779 nor n598 n827 ; n828
g780 nor a[22] n58 ; n829
g781 and a[9] n829_not ; n830
g782 and a[9]_not n829 ; n831
g783 nor n830 n831 ; n832
g784 nor n444 n832 ; n833
g785 and n828_not n833 ; n834
g786 and n828 n833_not ; n835
g787 nor n834 n835 ; n836
g788 and a[10] a[22] ; n837
g789 and a[10] n59_not ; n838
g790 and n666 n838_not ; n839
g791 nor n837 n839 ; n840
g792 nor n444 n840 ; n841
g793 and n836 n841 ; n842
g794 nor n834 n842 ; n843
g795 nor n695 n697 ; n844
g796 and n525_not n844 ; n845
g797 and n525 n700 ; n846
g798 and n665_not n695 ; n847
g799 and n529 n847 ; n848
g800 and n529_not n698 ; n849
g801 nor n848 n849 ; n850
g802 and n846_not n850 ; n851
g803 and n845_not n851 ; n852
g804 and n677_not n684 ; n853
g805 and n545 n677 ; n854
g806 and n669 n687 ; n855
g807 and n542 n669_not ; n856
g808 nor n855 n856 ; n857
g809 and n854_not n857 ; n858
g810 and n853_not n858 ; n859
g811 and n852 n859 ; n860
g812 and n786 n826_not ; n861
g813 and n786_not n826 ; n862
g814 nor n861 n862 ; n863
g815 and n786 n826 ; n864
g816 and n598 n864_not ; n865
g817 and n863 n865_not ; n866
g818 and n525_not n866 ; n867
g819 nor n828 n863 ; n868
g820 and n525 n828_not ; n869
g821 nor n868 n869 ; n870
g822 and n867_not n870 ; n871
g823 and n833_not n871 ; n872
g824 and n529_not n844 ; n873
g825 and n529 n700 ; n874
g826 and n677 n847 ; n875
g827 and n677_not n698 ; n876
g828 nor n875 n876 ; n877
g829 and n874_not n877 ; n878
g830 and n873_not n878 ; n879
g831 and n833 n871_not ; n880
g832 nor n872 n880 ; n881
g833 and n879 n881 ; n882
g834 nor n872 n882 ; n883
g835 nor n852 n859 ; n884
g836 nor n860 n884 ; n885
g837 and n883_not n885 ; n886
g838 nor n860 n886 ; n887
g839 nor n843 n887 ; n888
g840 nor n843 n888 ; n889
g841 nor n887 n888 ; n890
g842 nor n889 n890 ; n891
g843 nor n711 n713 ; n892
g844 nor n714 n892 ; n893
g845 and n891_not n893 ; n894
g846 nor n888 n894 ; n895
g847 nor n718 n720 ; n896
g848 nor n721 n896 ; n897
g849 and n895_not n897 ; n898
g850 and n669_not n684 ; n899
g851 and n545 n669 ; n900
g852 and n687 n840 ; n901
g853 and n542 n840_not ; n902
g854 nor n901 n902 ; n903
g855 and n900_not n903 ; n904
g856 and n899_not n904 ; n905
g857 nor n166 n446 ; n906
g858 and n145 n906 ; n907
g859 and n552_not n907 ; n908
g860 and n238_not n908 ; n909
g861 and n296_not n909 ; n910
g862 nor n174 n470 ; n911
g863 and n222_not n911 ; n912
g864 and n350_not n912 ; n913
g865 and n345_not n913 ; n914
g866 and n303 n914 ; n915
g867 and n323 n915 ; n916
g868 and n910 n916 ; n917
g869 and n152_not n917 ; n918
g870 and n196_not n918 ; n919
g871 and n186_not n919 ; n920
g872 and n504_not n920 ; n921
g873 and n495_not n921 ; n922
g874 and n154_not n922 ; n923
g875 nor n370 n468 ; n924
g876 and n347_not n924 ; n925
g877 and n445_not n925 ; n926
g878 and n127_not n407 ; n927
g879 and n216_not n927 ; n928
g880 and n589_not n928 ; n929
g881 and n367_not n929 ; n930
g882 nor n139 n327 ; n931
g883 and n562 n638 ; n932
g884 and n931 n932 ; n933
g885 and n930 n933 ; n934
g886 and n926 n934 ; n935
g887 and n219_not n935 ; n936
g888 and n299_not n936 ; n937
g889 and n148_not n937 ; n938
g890 nor n177 n214 ; n939
g891 and n218_not n939 ; n940
g892 and n192_not n940 ; n941
g893 and n133_not n941 ; n942
g894 and n736_not n942 ; n943
g895 and n342_not n943 ; n944
g896 nor n190 n394 ; n945
g897 and n235_not n945 ; n946
g898 nor n155 n405 ; n947
g899 and n351_not n947 ; n948
g900 and n496 n573 ; n949
g901 and n948 n949 ; n950
g902 and n946 n950 ; n951
g903 and n325 n951 ; n952
g904 and n944 n952 ; n953
g905 and n938 n953 ; n954
g906 and n923 n954 ; n955
g907 and n300_not n955 ; n956
g908 and n255_not n956 ; n957
g909 and n258_not n957 ; n958
g910 and n553_not n958 ; n959
g911 nor n169 n360 ; n960
g912 and n447_not n960 ; n961
g913 and n155_not n961 ; n962
g914 and n350_not n962 ; n963
g915 and n218_not n963 ; n964
g916 and n234_not n964 ; n965
g917 and n359_not n965 ; n966
g918 and n357_not n966 ; n967
g919 nor n133 n257 ; n968
g920 and n368_not n968 ; n969
g921 nor n469 n471 ; n970
g922 and n969 n970 ; n971
g923 and n144_not n971 ; n972
g924 and n327_not n972 ; n973
g925 and n446_not n973 ; n974
g926 and n315_not n974 ; n975
g927 nor n190 n302 ; n976
g928 and n174_not n976 ; n977
g929 and n191_not n977 ; n978
g930 and n168_not n978 ; n979
g931 nor n222 n408 ; n980
g932 and n394_not n980 ; n981
g933 and n228_not n981 ; n982
g934 and n417_not n982 ; n983
g935 nor n129 n178 ; n984
g936 and n196_not n984 ; n985
g937 and n449_not n985 ; n986
g938 and n256 n986 ; n987
g939 and n983 n987 ; n988
g940 and n926 n988 ; n989
g941 and n328_not n989 ; n990
g942 and n176_not n990 ; n991
g943 and n220_not n991 ; n992
g944 and n172_not n992 ; n993
g945 and n787 n993 ; n994
g946 and n223_not n994 ; n995
g947 and n337_not n995 ; n996
g948 and n175_not n996 ; n997
g949 and n552_not n997 ; n998
g950 and n351_not n998 ; n999
g951 and n979 n999 ; n1000
g952 and n141 n1000 ; n1001
g953 and n975 n1001 ; n1002
g954 and n967 n1002 ; n1003
g955 and n614 n1003 ; n1004
g956 and n299_not n1004 ; n1005
g957 and n503_not n1005 ; n1006
g958 and n367_not n1006 ; n1007
g959 nor n959 n1007 ; n1008
g960 nor n786 n1008 ; n1009
g961 nor a[22] n56 ; n1010
g962 and a[7] n1010_not ; n1011
g963 and a[7]_not n1010 ; n1012
g964 nor n1011 n1012 ; n1013
g965 nor n444 n1013 ; n1014
g966 and n1009_not n1014 ; n1015
g967 and n1009 n1014_not ; n1016
g968 nor n1015 n1016 ; n1017
g969 and a[8] a[22] ; n1018
g970 and a[8] n57_not ; n1019
g971 and n829 n1019_not ; n1020
g972 nor n1018 n1020 ; n1021
g973 and n1017 n1021_not ; n1022
g974 and n444_not n1022 ; n1023
g975 nor n1015 n1023 ; n1024
g976 and n905 n1024_not ; n1025
g977 and n684 n840_not ; n1026
g978 and n545 n840 ; n1027
g979 and n687 n832 ; n1028
g980 and n542 n832_not ; n1029
g981 nor n1028 n1029 ; n1030
g982 and n1027_not n1030 ; n1031
g983 and n1026_not n1031 ; n1032
g984 nor n863 n865 ; n1033
g985 and n525_not n1033 ; n1034
g986 and n525 n868 ; n1035
g987 and n828_not n863 ; n1036
g988 and n529 n1036 ; n1037
g989 and n529_not n866 ; n1038
g990 nor n1037 n1038 ; n1039
g991 and n1035_not n1039 ; n1040
g992 and n1034_not n1040 ; n1041
g993 and n677_not n844 ; n1042
g994 and n677 n700 ; n1043
g995 and n669 n847 ; n1044
g996 and n669_not n698 ; n1045
g997 nor n1044 n1045 ; n1046
g998 and n1043_not n1046 ; n1047
g999 and n1042_not n1047 ; n1048
g1000 and n1041 n1048_not ; n1049
g1001 and n1041_not n1048 ; n1050
g1002 nor n1049 n1050 ; n1051
g1003 and n1032 n1051_not ; n1052
g1004 and n1041 n1048 ; n1053
g1005 nor n1052 n1053 ; n1054
g1006 and n905 n1025_not ; n1055
g1007 nor n1024 n1025 ; n1056
g1008 nor n1055 n1056 ; n1057
g1009 nor n1054 n1057 ; n1058
g1010 nor n1025 n1058 ; n1059
g1011 nor n836 n841 ; n1060
g1012 nor n842 n1060 ; n1061
g1013 and n1059_not n1061 ; n1062
g1014 and n1059 n1061_not ; n1063
g1015 nor n1062 n1063 ; n1064
g1016 and n883 n885_not ; n1065
g1017 nor n886 n1065 ; n1066
g1018 and n1064 n1066 ; n1067
g1019 nor n1062 n1067 ; n1068
g1020 nor n891 n894 ; n1069
g1021 and n893 n894_not ; n1070
g1022 nor n1069 n1070 ; n1071
g1023 and n1068_not n1071 ; n1072
g1024 and n1068 n1071_not ; n1073
g1025 nor n1072 n1073 ; n1074
g1026 and n669_not n844 ; n1075
g1027 and n669 n700 ; n1076
g1028 and n840 n847 ; n1077
g1029 and n698 n840_not ; n1078
g1030 nor n1077 n1078 ; n1079
g1031 and n1076_not n1079 ; n1080
g1032 and n1075_not n1080 ; n1081
g1033 and n684 n832_not ; n1082
g1034 and n545 n832 ; n1083
g1035 and n687 n1021 ; n1084
g1036 and n542 n1021_not ; n1085
g1037 nor n1084 n1085 ; n1086
g1038 and n1083_not n1086 ; n1087
g1039 and n1082_not n1087 ; n1088
g1040 and n1081 n1088 ; n1089
g1041 nor n348 n495 ; n1090
g1042 and n335_not n1090 ; n1091
g1043 nor n226 n446 ; n1092
g1044 and n553_not n1092 ; n1093
g1045 nor n175 n343 ; n1094
g1046 and n503_not n1094 ; n1095
g1047 and n472_not n1095 ; n1096
g1048 and n1093 n1096 ; n1097
g1049 and n1091 n1097 ; n1098
g1050 and n983 n1098 ; n1099
g1051 and n149 n1099 ; n1100
g1052 and n196_not n1100 ; n1101
g1053 and n327_not n1101 ; n1102
g1054 and n212_not n1102 ; n1103
g1055 and n469_not n1103 ; n1104
g1056 and n118_not n395 ; n1105
g1057 and n235_not n1105 ; n1106
g1058 and n448 n1106 ; n1107
g1059 and n224_not n1107 ; n1108
g1060 and n460 n468_not ; n1109
g1061 and n176_not n1109 ; n1110
g1062 and n214_not n1110 ; n1111
g1063 and n218_not n1111 ; n1112
g1064 and n504_not n1112 ; n1113
g1065 and n358_not n1113 ; n1114
g1066 and n345_not n1114 ; n1115
g1067 nor n223 n599 ; n1116
g1068 nor n140 n336 ; n1117
g1069 and n1116 n1117 ; n1118
g1070 and n609 n1118 ; n1119
g1071 and n558 n1119 ; n1120
g1072 and n325 n1120 ; n1121
g1073 and n1115 n1121 ; n1122
g1074 and n1108 n1122 ; n1123
g1075 and n311 n1123 ; n1124
g1076 and n1104 n1124 ; n1125
g1077 and n188_not n1125 ; n1126
g1078 and n133_not n1126 ; n1127
g1079 and n206_not n1127 ; n1128
g1080 and n166_not n1128 ; n1129
g1081 and n552_not n1129 ; n1130
g1082 and n459 n1116 ; n1131
g1083 and n807 n1131 ; n1132
g1084 and n220_not n1132 ; n1133
g1085 and n394_not n1133 ; n1134
g1086 and n646 n948 ; n1135
g1087 and n314 n1135 ; n1136
g1088 and n1108 n1136 ; n1137
g1089 and n1134 n1137 ; n1138
g1090 and n129_not n1138 ; n1139
g1091 and n196_not n1139 ; n1140
g1092 and n150_not n1140 ; n1141
g1093 and n213_not n1141 ; n1142
g1094 and n169_not n1142 ; n1143
g1095 and n315_not n1143 ; n1144
g1096 and n326_not n1144 ; n1145
g1097 and n637 n911 ; n1146
g1098 and n194_not n1146 ; n1147
g1099 and n214_not n1147 ; n1148
g1100 and n348_not n1148 ; n1149
g1101 and n299_not n1149 ; n1150
g1102 and n552_not n1150 ; n1151
g1103 and n736_not n1151 ; n1152
g1104 and n560 n969 ; n1153
g1105 and n324_not n1153 ; n1154
g1106 and n1152 n1154 ; n1155
g1107 and n475 n1155 ; n1156
g1108 and n167_not n1156 ; n1157
g1109 and n336_not n1157 ; n1158
g1110 and n258_not n1158 ; n1159
g1111 and n345_not n1159 ; n1160
g1112 and n154_not n1160 ; n1161
g1113 and n215_not n1161 ; n1162
g1114 nor n208 n408 ; n1163
g1115 and n142_not n1163 ; n1164
g1116 and n111_not n1164 ; n1165
g1117 and n760 n1165 ; n1166
g1118 and n451 n1166 ; n1167
g1119 and n505 n1167 ; n1168
g1120 and n366 n1168 ; n1169
g1121 and n141 n1169 ; n1170
g1122 and n1162 n1170 ; n1171
g1123 and n1145 n1171 ; n1172
g1124 and n152_not n1172 ; n1173
g1125 and n219_not n1173 ; n1174
g1126 and n335_not n1174 ; n1175
g1127 nor n1130 n1175 ; n1176
g1128 nor n959 n1176 ; n1177
g1129 and n1130 n1177_not ; n1178
g1130 and n1130_not n1177 ; n1179
g1131 and a[6] a[22] ; n1180
g1132 and a[6] n55_not ; n1181
g1133 and n1010 n1181_not ; n1182
g1134 nor n1180 n1182 ; n1183
g1135 nor n444 n1183 ; n1184
g1136 and n1178_not n1184 ; n1185
g1137 and n1179_not n1185 ; n1186
g1138 nor n1178 n1186 ; n1187
g1139 nor n1081 n1088 ; n1188
g1140 nor n1089 n1188 ; n1189
g1141 and n1187_not n1189 ; n1190
g1142 nor n1089 n1190 ; n1191
g1143 and n959 n1007_not ; n1192
g1144 and n959_not n1007 ; n1193
g1145 nor n1192 n1193 ; n1194
g1146 and n959 n1007 ; n1195
g1147 and n786 n1195_not ; n1196
g1148 and n1194 n1196_not ; n1197
g1149 and n525_not n1197 ; n1198
g1150 nor n1009 n1194 ; n1199
g1151 and n525 n1009_not ; n1200
g1152 nor n1199 n1200 ; n1201
g1153 and n1198_not n1201 ; n1202
g1154 and n1014_not n1202 ; n1203
g1155 and n529_not n1033 ; n1204
g1156 and n529 n868 ; n1205
g1157 and n677 n1036 ; n1206
g1158 and n677_not n866 ; n1207
g1159 nor n1206 n1207 ; n1208
g1160 and n1205_not n1208 ; n1209
g1161 and n1204_not n1209 ; n1210
g1162 and n1014 n1202_not ; n1211
g1163 nor n1203 n1211 ; n1212
g1164 and n1210 n1212 ; n1213
g1165 nor n1203 n1213 ; n1214
g1166 nor n1191 n1214 ; n1215
g1167 nor n1191 n1215 ; n1216
g1168 nor n1214 n1215 ; n1217
g1169 nor n1216 n1217 ; n1218
g1170 nor n444 n1023 ; n1219
g1171 and n1021_not n1219 ; n1220
g1172 and n1017 n1023_not ; n1221
g1173 nor n1220 n1221 ; n1222
g1174 nor n1218 n1222 ; n1223
g1175 nor n1215 n1223 ; n1224
g1176 nor n879 n881 ; n1225
g1177 nor n882 n1225 ; n1226
g1178 and n1224_not n1226 ; n1227
g1179 nor n1054 n1058 ; n1228
g1180 nor n1057 n1058 ; n1229
g1181 nor n1228 n1229 ; n1230
g1182 and n1224 n1226_not ; n1231
g1183 nor n1227 n1231 ; n1232
g1184 and n1230_not n1232 ; n1233
g1185 nor n1227 n1233 ; n1234
g1186 nor n1064 n1066 ; n1235
g1187 nor n1067 n1235 ; n1236
g1188 and n1234_not n1236 ; n1237
g1189 and n1232 n1233_not ; n1238
g1190 nor n1230 n1233 ; n1239
g1191 nor n1238 n1239 ; n1240
g1192 nor n1194 n1196 ; n1241
g1193 and n525_not n1241 ; n1242
g1194 and n525 n1199 ; n1243
g1195 and n1009_not n1194 ; n1244
g1196 and n529 n1244 ; n1245
g1197 and n529_not n1197 ; n1246
g1198 nor n1245 n1246 ; n1247
g1199 and n1243_not n1247 ; n1248
g1200 and n1242_not n1248 ; n1249
g1201 and n840_not n844 ; n1250
g1202 and n700 n840 ; n1251
g1203 and n832 n847 ; n1252
g1204 and n698 n832_not ; n1253
g1205 nor n1252 n1253 ; n1254
g1206 and n1251_not n1254 ; n1255
g1207 and n1250_not n1255 ; n1256
g1208 and n684 n1021_not ; n1257
g1209 and n545 n1021 ; n1258
g1210 and n687 n1013 ; n1259
g1211 and n542 n1013_not ; n1260
g1212 nor n1259 n1260 ; n1261
g1213 and n1258_not n1261 ; n1262
g1214 and n1257_not n1262 ; n1263
g1215 and n1256 n1263_not ; n1264
g1216 and n1256_not n1263 ; n1265
g1217 nor n1264 n1265 ; n1266
g1218 and n1249 n1266_not ; n1267
g1219 and n1256 n1263 ; n1268
g1220 nor n1267 n1268 ; n1269
g1221 nor n1210 n1212 ; n1270
g1222 nor n1213 n1270 ; n1271
g1223 and n1269_not n1271 ; n1272
g1224 nor n1269 n1272 ; n1273
g1225 and n1271 n1272_not ; n1274
g1226 nor n1273 n1274 ; n1275
g1227 and n1187 n1189_not ; n1276
g1228 nor n1190 n1276 ; n1277
g1229 and n1275_not n1277 ; n1278
g1230 nor n1272 n1278 ; n1279
g1231 and n1032 n1052_not ; n1280
g1232 nor n1051 n1052 ; n1281
g1233 nor n1280 n1281 ; n1282
g1234 nor n1279 n1282 ; n1283
g1235 nor n1279 n1283 ; n1284
g1236 nor n1282 n1283 ; n1285
g1237 nor n1284 n1285 ; n1286
g1238 nor n1218 n1223 ; n1287
g1239 nor n1222 n1223 ; n1288
g1240 nor n1287 n1288 ; n1289
g1241 nor n1286 n1289 ; n1290
g1242 nor n1283 n1290 ; n1291
g1243 nor n1240 n1291 ; n1292
g1244 nor n1240 n1292 ; n1293
g1245 nor n1291 n1292 ; n1294
g1246 nor n1293 n1294 ; n1295
g1247 and n677_not n1033 ; n1296
g1248 and n677 n868 ; n1297
g1249 and n669 n1036 ; n1298
g1250 and n669_not n866 ; n1299
g1251 nor n1298 n1299 ; n1300
g1252 and n1297_not n1300 ; n1301
g1253 and n1296_not n1301 ; n1302
g1254 and n1179_not n1187 ; n1303
g1255 and n1184 n1186_not ; n1304
g1256 nor n1303 n1304 ; n1305
g1257 and n1302 n1305_not ; n1306
g1258 nor n275 n444 ; n1307
g1259 and n1130_not n1307 ; n1308
g1260 and n1130 n1307_not ; n1309
g1261 and n1130 n1175_not ; n1310
g1262 and n1130_not n1175 ; n1311
g1263 nor n1310 n1311 ; n1312
g1264 and n1130 n1175 ; n1313
g1265 and n959 n1313_not ; n1314
g1266 and n1312 n1314_not ; n1315
g1267 and n525_not n1315 ; n1316
g1268 nor n1177 n1312 ; n1317
g1269 and n525 n1177_not ; n1318
g1270 nor n1317 n1318 ; n1319
g1271 and n1316_not n1319 ; n1320
g1272 and n1308_not n1320 ; n1321
g1273 and n1309_not n1321 ; n1322
g1274 nor n1308 n1322 ; n1323
g1275 and n1302_not n1305 ; n1324
g1276 nor n1306 n1324 ; n1325
g1277 and n1323_not n1325 ; n1326
g1278 nor n1306 n1326 ; n1327
g1279 and n529_not n1241 ; n1328
g1280 and n529 n1199 ; n1329
g1281 and n677 n1244 ; n1330
g1282 and n677_not n1197 ; n1331
g1283 nor n1330 n1331 ; n1332
g1284 and n1329_not n1332 ; n1333
g1285 and n1328_not n1333 ; n1334
g1286 and n669_not n1033 ; n1335
g1287 and n669 n868 ; n1336
g1288 and n840 n1036 ; n1337
g1289 and n840_not n866 ; n1338
g1290 nor n1337 n1338 ; n1339
g1291 and n1336_not n1339 ; n1340
g1292 and n1335_not n1340 ; n1341
g1293 and n1334 n1341 ; n1342
g1294 and n832_not n844 ; n1343
g1295 and n700 n832 ; n1344
g1296 and n847 n1021 ; n1345
g1297 and n698 n1021_not ; n1346
g1298 nor n1345 n1346 ; n1347
g1299 and n1344_not n1347 ; n1348
g1300 and n1343_not n1348 ; n1349
g1301 and n1334 n1341_not ; n1350
g1302 and n1334_not n1341 ; n1351
g1303 nor n1350 n1351 ; n1352
g1304 and n1349 n1352_not ; n1353
g1305 nor n1342 n1353 ; n1354
g1306 and n1249_not n1266 ; n1355
g1307 nor n1267 n1355 ; n1356
g1308 and n1354_not n1356 ; n1357
g1309 and n684 n1013_not ; n1358
g1310 and n545 n1013 ; n1359
g1311 and n687 n1183 ; n1360
g1312 and n542 n1183_not ; n1361
g1313 nor n1360 n1361 ; n1362
g1314 and n1359_not n1362 ; n1363
g1315 and n1358_not n1363 ; n1364
g1316 nor n279 n444 ; n1365
g1317 and n1130_not n1365 ; n1366
g1318 and n1130 n1365_not ; n1367
g1319 nor n1312 n1314 ; n1368
g1320 and n525_not n1368 ; n1369
g1321 and n525 n1317 ; n1370
g1322 and n1177_not n1312 ; n1371
g1323 and n529 n1371 ; n1372
g1324 and n529_not n1315 ; n1373
g1325 nor n1372 n1373 ; n1374
g1326 and n1370_not n1374 ; n1375
g1327 and n1369_not n1375 ; n1376
g1328 and n1366_not n1376 ; n1377
g1329 and n1367_not n1377 ; n1378
g1330 nor n1366 n1378 ; n1379
g1331 and n1364 n1379_not ; n1380
g1332 and n1364_not n1379 ; n1381
g1333 nor n1380 n1381 ; n1382
g1334 and n840_not n1033 ; n1383
g1335 and n840 n868 ; n1384
g1336 and n832 n1036 ; n1385
g1337 and n832_not n866 ; n1386
g1338 nor n1385 n1386 ; n1387
g1339 and n1384_not n1387 ; n1388
g1340 and n1383_not n1388 ; n1389
g1341 and n677_not n1241 ; n1390
g1342 and n677 n1199 ; n1391
g1343 and n669 n1244 ; n1392
g1344 and n669_not n1197 ; n1393
g1345 nor n1392 n1393 ; n1394
g1346 and n1391_not n1394 ; n1395
g1347 and n1390_not n1395 ; n1396
g1348 and n1389 n1396 ; n1397
g1349 and n844 n1021_not ; n1398
g1350 and n700 n1021 ; n1399
g1351 and n847 n1013 ; n1400
g1352 and n698 n1013_not ; n1401
g1353 nor n1400 n1401 ; n1402
g1354 and n1399_not n1402 ; n1403
g1355 and n1398_not n1403 ; n1404
g1356 and n1389_not n1396 ; n1405
g1357 and n1389 n1396_not ; n1406
g1358 nor n1405 n1406 ; n1407
g1359 and n1404 n1407_not ; n1408
g1360 nor n1397 n1408 ; n1409
g1361 and n1382 n1409_not ; n1410
g1362 nor n1380 n1410 ; n1411
g1363 and n1354 n1356_not ; n1412
g1364 nor n1357 n1412 ; n1413
g1365 and n1411_not n1413 ; n1414
g1366 nor n1357 n1414 ; n1415
g1367 nor n1327 n1415 ; n1416
g1368 nor n1327 n1416 ; n1417
g1369 nor n1415 n1416 ; n1418
g1370 nor n1417 n1418 ; n1419
g1371 and n1277 n1278_not ; n1420
g1372 nor n1275 n1278 ; n1421
g1373 nor n1420 n1421 ; n1422
g1374 nor n1419 n1422 ; n1423
g1375 nor n1416 n1423 ; n1424
g1376 and n1286_not n1289 ; n1425
g1377 and n1286 n1289_not ; n1426
g1378 nor n1425 n1426 ; n1427
g1379 nor n1424 n1427 ; n1428
g1380 nor n1419 n1423 ; n1429
g1381 nor n1422 n1423 ; n1430
g1382 nor n1429 n1430 ; n1431
g1383 and n1309_not n1323 ; n1432
g1384 and n1320 n1322_not ; n1433
g1385 nor n1432 n1433 ; n1434
g1386 and n1349 n1353_not ; n1435
g1387 nor n1352 n1353 ; n1436
g1388 nor n1435 n1436 ; n1437
g1389 nor n1434 n1437 ; n1438
g1390 nor n1434 n1438 ; n1439
g1391 nor n1437 n1438 ; n1440
g1392 nor n1439 n1440 ; n1441
g1393 and n684 n1183_not ; n1442
g1394 and n545 n1183 ; n1443
g1395 and n275 n687 ; n1444
g1396 and n275_not n542 ; n1445
g1397 nor n1444 n1445 ; n1446
g1398 and n1443_not n1446 ; n1447
g1399 and n1442_not n1447 ; n1448
g1400 nor n286 n444 ; n1449
g1401 and n221_not n809 ; n1450
g1402 and n174_not n1450 ; n1451
g1403 and n300_not n1451 ; n1452
g1404 and n123_not n1452 ; n1453
g1405 and n212_not n1453 ; n1454
g1406 and n347_not n1454 ; n1455
g1407 and n552_not n1455 ; n1456
g1408 and n553_not n1456 ; n1457
g1409 nor n220 n350 ; n1458
g1410 and n315_not n1458 ; n1459
g1411 and n432 n584 ; n1460
g1412 and n1459 n1460 ; n1461
g1413 and n968 n1461 ; n1462
g1414 and n644 n1462 ; n1463
g1415 and n337_not n1463 ; n1464
g1416 and n214_not n1464 ; n1465
g1417 and n417_not n1465 ; n1466
g1418 and n234_not n1466 ; n1467
g1419 and n367_not n1467 ; n1468
g1420 nor n324 n360 ; n1469
g1421 and n446_not n1469 ; n1470
g1422 and n172_not n1470 ; n1471
g1423 and n503_not n1471 ; n1472
g1424 and n356_not n1472 ; n1473
g1425 and n216_not n1473 ; n1474
g1426 and n342_not n1474 ; n1475
g1427 and n154_not n1475 ; n1476
g1428 and n373 n1476 ; n1477
g1429 and n1468 n1477 ; n1478
g1430 and n421 n1478 ; n1479
g1431 and n1457 n1479 ; n1480
g1432 and n178_not n1480 ; n1481
g1433 and n208_not n1481 ; n1482
g1434 and n118_not n1482 ; n1483
g1435 and n361_not n1483 ; n1484
g1436 and n258_not n1484 ; n1485
g1437 and n599_not n1485 ; n1486
g1438 and n211_not n1486 ; n1487
g1439 and n525_not n1487 ; n1488
g1440 nor n1130 n1488 ; n1489
g1441 and n1449 n1489 ; n1490
g1442 and n529_not n1368 ; n1491
g1443 and n529 n1317 ; n1492
g1444 and n677 n1371 ; n1493
g1445 and n677_not n1315 ; n1494
g1446 nor n1493 n1494 ; n1495
g1447 and n1492_not n1495 ; n1496
g1448 and n1491_not n1496 ; n1497
g1449 nor n1449 n1489 ; n1498
g1450 nor n1490 n1498 ; n1499
g1451 and n1497 n1499 ; n1500
g1452 nor n1490 n1500 ; n1501
g1453 and n1448 n1501_not ; n1502
g1454 and n1448_not n1501 ; n1503
g1455 nor n1502 n1503 ; n1504
g1456 and n832_not n1033 ; n1505
g1457 and n832 n868 ; n1506
g1458 and n1021 n1036 ; n1507
g1459 and n866 n1021_not ; n1508
g1460 nor n1507 n1508 ; n1509
g1461 and n1506_not n1509 ; n1510
g1462 and n1505_not n1510 ; n1511
g1463 and n669_not n1241 ; n1512
g1464 and n669 n1199 ; n1513
g1465 and n840 n1244 ; n1514
g1466 and n840_not n1197 ; n1515
g1467 nor n1514 n1515 ; n1516
g1468 and n1513_not n1516 ; n1517
g1469 and n1512_not n1517 ; n1518
g1470 and n1511 n1518 ; n1519
g1471 and n844 n1013_not ; n1520
g1472 and n700 n1013 ; n1521
g1473 and n847 n1183 ; n1522
g1474 and n698 n1183_not ; n1523
g1475 nor n1522 n1523 ; n1524
g1476 and n1521_not n1524 ; n1525
g1477 and n1520_not n1525 ; n1526
g1478 and n1511_not n1518 ; n1527
g1479 and n1511 n1518_not ; n1528
g1480 nor n1527 n1528 ; n1529
g1481 and n1526 n1529_not ; n1530
g1482 nor n1519 n1530 ; n1531
g1483 and n1504 n1531_not ; n1532
g1484 nor n1502 n1532 ; n1533
g1485 nor n1441 n1533 ; n1534
g1486 nor n1438 n1534 ; n1535
g1487 and n1323 n1325_not ; n1536
g1488 nor n1326 n1536 ; n1537
g1489 and n1535_not n1537 ; n1538
g1490 and n1535 n1537_not ; n1539
g1491 nor n1538 n1539 ; n1540
g1492 and n1411 n1413_not ; n1541
g1493 nor n1414 n1541 ; n1542
g1494 and n1540 n1542 ; n1543
g1495 nor n1538 n1543 ; n1544
g1496 nor n1431 n1544 ; n1545
g1497 and n1431 n1544_not ; n1546
g1498 and n1431_not n1544 ; n1547
g1499 nor n1546 n1547 ; n1548
g1500 and n1130 n1487_not ; n1549
g1501 nor n1487 n1549 ; n1550
g1502 and n525_not n1550 ; n1551
g1503 and n525 n1549 ; n1552
g1504 and n529 n1130_not ; n1553
g1505 and n1487 n1553_not ; n1554
g1506 nor n1552 n1554 ; n1555
g1507 and n1551_not n1555 ; n1556
g1508 and n286_not n684 ; n1557
g1509 and n286 n544_not ; n1558
g1510 nor n687 n1558 ; n1559
g1511 and n1557_not n1559 ; n1560
g1512 and n544 n1560 ; n1561
g1513 and n1556 n1561 ; n1562
g1514 and n275_not n684 ; n1563
g1515 and n275 n545 ; n1564
g1516 and n279 n687 ; n1565
g1517 and n279_not n542 ; n1566
g1518 nor n1565 n1566 ; n1567
g1519 and n1564_not n1567 ; n1568
g1520 and n1563_not n1568 ; n1569
g1521 and n1562 n1569 ; n1570
g1522 and n840_not n1241 ; n1571
g1523 and n840 n1199 ; n1572
g1524 and n832 n1244 ; n1573
g1525 and n832_not n1197 ; n1574
g1526 nor n1573 n1574 ; n1575
g1527 and n1572_not n1575 ; n1576
g1528 and n1571_not n1576 ; n1577
g1529 and n1021_not n1033 ; n1578
g1530 and n868 n1021 ; n1579
g1531 and n1013 n1036 ; n1580
g1532 and n866 n1013_not ; n1581
g1533 nor n1580 n1581 ; n1582
g1534 and n1579_not n1582 ; n1583
g1535 and n1578_not n1583 ; n1584
g1536 and n844 n1183_not ; n1585
g1537 and n700 n1183 ; n1586
g1538 and n275 n847 ; n1587
g1539 and n275_not n698 ; n1588
g1540 nor n1587 n1588 ; n1589
g1541 and n1586_not n1589 ; n1590
g1542 and n1585_not n1590 ; n1591
g1543 and n1584 n1591_not ; n1592
g1544 and n1584_not n1591 ; n1593
g1545 nor n1592 n1593 ; n1594
g1546 and n1577 n1594_not ; n1595
g1547 and n1584 n1591 ; n1596
g1548 nor n1595 n1596 ; n1597
g1549 nor n1562 n1569 ; n1598
g1550 nor n1570 n1598 ; n1599
g1551 and n1597_not n1599 ; n1600
g1552 nor n1570 n1600 ; n1601
g1553 and n1367_not n1379 ; n1602
g1554 and n1376 n1378_not ; n1603
g1555 nor n1602 n1603 ; n1604
g1556 and n1601 n1604_not ; n1605
g1557 and n1601_not n1604 ; n1606
g1558 nor n1605 n1606 ; n1607
g1559 and n1404 n1408_not ; n1608
g1560 nor n1407 n1408 ; n1609
g1561 nor n1608 n1609 ; n1610
g1562 nor n1607 n1610 ; n1611
g1563 nor n1601 n1604 ; n1612
g1564 nor n1611 n1612 ; n1613
g1565 and n1382_not n1409 ; n1614
g1566 nor n1410 n1614 ; n1615
g1567 and n1613_not n1615 ; n1616
g1568 and n1441 n1533_not ; n1617
g1569 and n1441_not n1533 ; n1618
g1570 nor n1617 n1618 ; n1619
g1571 and n1613 n1615_not ; n1620
g1572 nor n1616 n1620 ; n1621
g1573 and n1619_not n1621 ; n1622
g1574 nor n1616 n1622 ; n1623
g1575 nor n1540 n1542 ; n1624
g1576 nor n1543 n1624 ; n1625
g1577 and n1623_not n1625 ; n1626
g1578 and n677_not n1368 ; n1627
g1579 and n677 n1317 ; n1628
g1580 and n669 n1371 ; n1629
g1581 and n669_not n1315 ; n1630
g1582 nor n1629 n1630 ; n1631
g1583 and n1628_not n1631 ; n1632
g1584 and n1627_not n1632 ; n1633
g1585 and n279_not n684 ; n1634
g1586 and n279 n545 ; n1635
g1587 and n286 n687 ; n1636
g1588 and n286_not n542 ; n1637
g1589 nor n1636 n1637 ; n1638
g1590 and n1635_not n1638 ; n1639
g1591 and n1634_not n1639 ; n1640
g1592 and n1633 n1640 ; n1641
g1593 nor n1556 n1561 ; n1642
g1594 nor n1562 n1642 ; n1643
g1595 nor n1633 n1640 ; n1644
g1596 nor n1641 n1644 ; n1645
g1597 and n1643 n1645 ; n1646
g1598 nor n1641 n1646 ; n1647
g1599 nor n1497 n1499 ; n1648
g1600 nor n1500 n1648 ; n1649
g1601 and n1647_not n1649 ; n1650
g1602 and n1647 n1649_not ; n1651
g1603 nor n1650 n1651 ; n1652
g1604 and n1526 n1530_not ; n1653
g1605 nor n1529 n1530 ; n1654
g1606 nor n1653 n1654 ; n1655
g1607 and n1652 n1655_not ; n1656
g1608 nor n1650 n1656 ; n1657
g1609 and n1504_not n1531 ; n1658
g1610 nor n1532 n1658 ; n1659
g1611 and n1657_not n1659 ; n1660
g1612 and n1657 n1659_not ; n1661
g1613 nor n1660 n1661 ; n1662
g1614 and n1607 n1610 ; n1663
g1615 nor n1611 n1663 ; n1664
g1616 and n1662 n1664 ; n1665
g1617 nor n1660 n1665 ; n1666
g1618 and n1619 n1621_not ; n1667
g1619 nor n1622 n1667 ; n1668
g1620 and n1666_not n1668 ; n1669
g1621 and n677_not n1550 ; n1670
g1622 and n677 n1549 ; n1671
g1623 and n669 n1130_not ; n1672
g1624 and n1487 n1672_not ; n1673
g1625 nor n1671 n1673 ; n1674
g1626 and n1670_not n1674 ; n1675
g1627 and n286_not n844 ; n1676
g1628 and n286 n665_not ; n1677
g1629 nor n847 n1677 ; n1678
g1630 and n1676_not n1678 ; n1679
g1631 and n665 n1679 ; n1680
g1632 and n1675 n1680 ; n1681
g1633 and n832_not n1241 ; n1682
g1634 and n832 n1199 ; n1683
g1635 and n1021 n1244 ; n1684
g1636 and n1021_not n1197 ; n1685
g1637 nor n1684 n1685 ; n1686
g1638 and n1683_not n1686 ; n1687
g1639 and n1682_not n1687 ; n1688
g1640 and n1013_not n1033 ; n1689
g1641 and n868 n1013 ; n1690
g1642 and n1036 n1183 ; n1691
g1643 and n866 n1183_not ; n1692
g1644 nor n1691 n1692 ; n1693
g1645 and n1690_not n1693 ; n1694
g1646 and n1689_not n1694 ; n1695
g1647 and n1688 n1695_not ; n1696
g1648 and n1688_not n1695 ; n1697
g1649 nor n1696 n1697 ; n1698
g1650 and n1681 n1698_not ; n1699
g1651 and n1688 n1695 ; n1700
g1652 nor n1699 n1700 ; n1701
g1653 and n275_not n844 ; n1702
g1654 and n275 n700 ; n1703
g1655 and n279 n847 ; n1704
g1656 and n279_not n698 ; n1705
g1657 nor n1704 n1705 ; n1706
g1658 and n1703_not n1706 ; n1707
g1659 and n1702_not n1707 ; n1708
g1660 and n529_not n1550 ; n1709
g1661 and n529 n1549 ; n1710
g1662 and n677 n1130_not ; n1711
g1663 and n1487 n1711_not ; n1712
g1664 nor n1710 n1712 ; n1713
g1665 and n1709_not n1713 ; n1714
g1666 and n669_not n1368 ; n1715
g1667 and n669 n1317 ; n1716
g1668 and n840 n1371 ; n1717
g1669 and n840_not n1315 ; n1718
g1670 nor n1717 n1718 ; n1719
g1671 and n1716_not n1719 ; n1720
g1672 and n1715_not n1720 ; n1721
g1673 and n1714 n1721_not ; n1722
g1674 and n1714_not n1721 ; n1723
g1675 nor n1722 n1723 ; n1724
g1676 and n1708 n1724_not ; n1725
g1677 and n1714 n1721 ; n1726
g1678 nor n1725 n1726 ; n1727
g1679 nor n1701 n1727 ; n1728
g1680 nor n1701 n1728 ; n1729
g1681 nor n1727 n1728 ; n1730
g1682 nor n1729 n1730 ; n1731
g1683 and n1577 n1595_not ; n1732
g1684 nor n1594 n1595 ; n1733
g1685 nor n1732 n1733 ; n1734
g1686 nor n1731 n1734 ; n1735
g1687 nor n1728 n1735 ; n1736
g1688 and n1597 n1599_not ; n1737
g1689 nor n1600 n1737 ; n1738
g1690 and n1736_not n1738 ; n1739
g1691 and n1652 n1656_not ; n1740
g1692 nor n1655 n1656 ; n1741
g1693 nor n1740 n1741 ; n1742
g1694 and n1736 n1738_not ; n1743
g1695 nor n1739 n1743 ; n1744
g1696 and n1742_not n1744 ; n1745
g1697 nor n1739 n1745 ; n1746
g1698 nor n1662 n1664 ; n1747
g1699 nor n1665 n1747 ; n1748
g1700 and n1746_not n1748 ; n1749
g1701 nor n544 n1560 ; n1750
g1702 and n1021_not n1241 ; n1751
g1703 and n1021 n1199 ; n1752
g1704 and n1013 n1244 ; n1753
g1705 and n1013_not n1197 ; n1754
g1706 nor n1753 n1754 ; n1755
g1707 and n1752_not n1755 ; n1756
g1708 and n1751_not n1756 ; n1757
g1709 and n840_not n1368 ; n1758
g1710 and n840 n1317 ; n1759
g1711 and n832 n1371 ; n1760
g1712 and n832_not n1315 ; n1761
g1713 nor n1760 n1761 ; n1762
g1714 and n1759_not n1762 ; n1763
g1715 and n1758_not n1763 ; n1764
g1716 and n1033 n1183_not ; n1765
g1717 and n868 n1183 ; n1766
g1718 and n275 n1036 ; n1767
g1719 and n275_not n866 ; n1768
g1720 nor n1767 n1768 ; n1769
g1721 and n1766_not n1769 ; n1770
g1722 and n1765_not n1770 ; n1771
g1723 and n1764 n1771_not ; n1772
g1724 and n1764_not n1771 ; n1773
g1725 nor n1772 n1773 ; n1774
g1726 and n1757 n1774_not ; n1775
g1727 and n1764 n1771 ; n1776
g1728 nor n1775 n1776 ; n1777
g1729 nor n1561 n1777 ; n1778
g1730 and n1750_not n1778 ; n1779
g1731 nor n1561 n1779 ; n1780
g1732 and n1750_not n1780 ; n1781
g1733 nor n1777 n1779 ; n1782
g1734 nor n1781 n1782 ; n1783
g1735 and n1681_not n1698 ; n1784
g1736 nor n1699 n1784 ; n1785
g1737 and n1783_not n1785 ; n1786
g1738 nor n1779 n1786 ; n1787
g1739 and n1643 n1646_not ; n1788
g1740 and n1644_not n1647 ; n1789
g1741 nor n1788 n1789 ; n1790
g1742 and n1787_not n1790 ; n1791
g1743 and n1787 n1790_not ; n1792
g1744 nor n1791 n1792 ; n1793
g1745 nor n1731 n1735 ; n1794
g1746 nor n1734 n1735 ; n1795
g1747 nor n1794 n1795 ; n1796
g1748 nor n1793 n1796 ; n1797
g1749 nor n1787 n1790 ; n1798
g1750 nor n1797 n1798 ; n1799
g1751 and n1742 n1744_not ; n1800
g1752 nor n1745 n1800 ; n1801
g1753 and n1799_not n1801 ; n1802
g1754 and n669_not n1550 ; n1803
g1755 and n669 n1549 ; n1804
g1756 and n840 n1130_not ; n1805
g1757 and n1487 n1805_not ; n1806
g1758 nor n1804 n1806 ; n1807
g1759 and n1803_not n1807 ; n1808
g1760 and n832_not n1368 ; n1809
g1761 and n832 n1317 ; n1810
g1762 and n1021 n1371 ; n1811
g1763 and n1021_not n1315 ; n1812
g1764 nor n1811 n1812 ; n1813
g1765 and n1810_not n1813 ; n1814
g1766 and n1809_not n1814 ; n1815
g1767 and n1808 n1815 ; n1816
g1768 and n1013_not n1241 ; n1817
g1769 and n1013 n1199 ; n1818
g1770 and n1183 n1244 ; n1819
g1771 and n1183_not n1197 ; n1820
g1772 nor n1819 n1820 ; n1821
g1773 and n1818_not n1821 ; n1822
g1774 and n1817_not n1822 ; n1823
g1775 and n1808 n1815_not ; n1824
g1776 and n1808_not n1815 ; n1825
g1777 nor n1824 n1825 ; n1826
g1778 and n1823 n1826_not ; n1827
g1779 nor n1816 n1827 ; n1828
g1780 and n279_not n844 ; n1829
g1781 and n279 n700 ; n1830
g1782 and n286 n847 ; n1831
g1783 and n286_not n698 ; n1832
g1784 nor n1831 n1832 ; n1833
g1785 and n1830_not n1833 ; n1834
g1786 and n1829_not n1834 ; n1835
g1787 nor n1675 n1680 ; n1836
g1788 nor n1681 n1836 ; n1837
g1789 and n1835 n1837_not ; n1838
g1790 and n1835_not n1837 ; n1839
g1791 nor n1838 n1839 ; n1840
g1792 nor n1828 n1840 ; n1841
g1793 and n1835 n1837 ; n1842
g1794 nor n1841 n1842 ; n1843
g1795 and n1708 n1725_not ; n1844
g1796 nor n1724 n1725 ; n1845
g1797 nor n1844 n1845 ; n1846
g1798 nor n1843 n1846 ; n1847
g1799 nor n1783 n1786 ; n1848
g1800 and n1785 n1786_not ; n1849
g1801 nor n1848 n1849 ; n1850
g1802 nor n1843 n1847 ; n1851
g1803 nor n1846 n1847 ; n1852
g1804 nor n1851 n1852 ; n1853
g1805 nor n1850 n1853 ; n1854
g1806 nor n1847 n1854 ; n1855
g1807 and n275_not n1033 ; n1856
g1808 and n275 n868 ; n1857
g1809 and n279 n1036 ; n1858
g1810 and n279_not n866 ; n1859
g1811 nor n1858 n1859 ; n1860
g1812 and n1857_not n1860 ; n1861
g1813 and n1856_not n1861 ; n1862
g1814 and n840_not n1550 ; n1863
g1815 and n840 n1549 ; n1864
g1816 and n832 n1130_not ; n1865
g1817 and n1487 n1865_not ; n1866
g1818 nor n1864 n1866 ; n1867
g1819 and n1863_not n1867 ; n1868
g1820 and n286_not n1033 ; n1869
g1821 and n286 n828_not ; n1870
g1822 nor n1036 n1870 ; n1871
g1823 and n1869_not n1871 ; n1872
g1824 and n828 n1872 ; n1873
g1825 and n1868 n1873 ; n1874
g1826 and n1862 n1874 ; n1875
g1827 and n1862_not n1874 ; n1876
g1828 and n1862 n1874_not ; n1877
g1829 nor n1876 n1877 ; n1878
g1830 nor n286 n695 ; n1879
g1831 and n1878_not n1879 ; n1880
g1832 nor n1875 n1880 ; n1881
g1833 and n1757_not n1774 ; n1882
g1834 nor n1775 n1882 ; n1883
g1835 and n1881_not n1883 ; n1884
g1836 and n1881 n1883_not ; n1885
g1837 nor n1884 n1885 ; n1886
g1838 and n1828 n1840 ; n1887
g1839 nor n1841 n1887 ; n1888
g1840 nor n1886 n1888 ; n1889
g1841 and n1886 n1888 ; n1890
g1842 and n279_not n1033 ; n1891
g1843 and n279 n868 ; n1892
g1844 and n286 n1036 ; n1893
g1845 and n286_not n866 ; n1894
g1846 nor n1893 n1894 ; n1895
g1847 and n1892_not n1895 ; n1896
g1848 and n1891_not n1896 ; n1897
g1849 and n1021_not n1368 ; n1898
g1850 and n1021 n1317 ; n1899
g1851 and n1013 n1371 ; n1900
g1852 and n1013_not n1315 ; n1901
g1853 nor n1900 n1901 ; n1902
g1854 and n1899_not n1902 ; n1903
g1855 and n1898_not n1903 ; n1904
g1856 and n1183_not n1241 ; n1905
g1857 and n1183 n1199 ; n1906
g1858 and n275 n1244 ; n1907
g1859 and n275_not n1197 ; n1908
g1860 nor n1907 n1908 ; n1909
g1861 and n1906_not n1909 ; n1910
g1862 and n1905_not n1910 ; n1911
g1863 and n1904 n1911_not ; n1912
g1864 and n1904_not n1911 ; n1913
g1865 nor n1912 n1913 ; n1914
g1866 and n1897 n1914_not ; n1915
g1867 and n1904 n1911 ; n1916
g1868 nor n1915 n1916 ; n1917
g1869 and n1823_not n1826 ; n1918
g1870 nor n1827 n1918 ; n1919
g1871 and n1917_not n1919 ; n1920
g1872 and n1878 n1879_not ; n1921
g1873 nor n1880 n1921 ; n1922
g1874 nor n1917 n1920 ; n1923
g1875 and n1919 n1920_not ; n1924
g1876 nor n1923 n1924 ; n1925
g1877 and n1922 n1925_not ; n1926
g1878 nor n1920 n1926 ; n1927
g1879 nor n828 n1872 ; n1928
g1880 and n1021_not n1550 ; n1929
g1881 and n1021 n1549 ; n1930
g1882 and n1013 n1130_not ; n1931
g1883 and n1487 n1931_not ; n1932
g1884 nor n1930 n1932 ; n1933
g1885 and n1929_not n1933 ; n1934
g1886 and n286_not n1241 ; n1935
g1887 and n286 n1009_not ; n1936
g1888 nor n1244 n1936 ; n1937
g1889 and n1935_not n1937 ; n1938
g1890 and n1009 n1938 ; n1939
g1891 and n1934 n1939 ; n1940
g1892 and n1873_not n1940 ; n1941
g1893 and n1928_not n1941 ; n1942
g1894 and n1183_not n1368 ; n1943
g1895 and n1183 n1317 ; n1944
g1896 and n275 n1371 ; n1945
g1897 and n275_not n1315 ; n1946
g1898 nor n1945 n1946 ; n1947
g1899 and n1944_not n1947 ; n1948
g1900 and n1943_not n1948 ; n1949
g1901 and n279_not n1241 ; n1950
g1902 and n279 n1199 ; n1951
g1903 and n286 n1244 ; n1952
g1904 and n286_not n1197 ; n1953
g1905 nor n1952 n1953 ; n1954
g1906 and n1951_not n1954 ; n1955
g1907 and n1950_not n1955 ; n1956
g1908 and n1949 n1956 ; n1957
g1909 nor n1934 n1939 ; n1958
g1910 nor n1940 n1958 ; n1959
g1911 nor n1949 n1956 ; n1960
g1912 nor n1957 n1960 ; n1961
g1913 and n1959 n1961 ; n1962
g1914 nor n1957 n1962 ; n1963
g1915 and n1940 n1942_not ; n1964
g1916 nor n1873 n1942 ; n1965
g1917 and n1928_not n1965 ; n1966
g1918 nor n1964 n1966 ; n1967
g1919 nor n1963 n1967 ; n1968
g1920 nor n1942 n1968 ; n1969
g1921 and n275_not n1241 ; n1970
g1922 and n275 n1199 ; n1971
g1923 and n279 n1244 ; n1972
g1924 and n279_not n1197 ; n1973
g1925 nor n1972 n1973 ; n1974
g1926 and n1971_not n1974 ; n1975
g1927 and n1970_not n1975 ; n1976
g1928 and n1013_not n1368 ; n1977
g1929 and n1013 n1317 ; n1978
g1930 and n1183 n1371 ; n1979
g1931 and n1183_not n1315 ; n1980
g1932 nor n1979 n1980 ; n1981
g1933 and n1978_not n1981 ; n1982
g1934 and n1977_not n1982 ; n1983
g1935 and n832_not n1550 ; n1984
g1936 and n832 n1549 ; n1985
g1937 and n1021 n1130_not ; n1986
g1938 and n1487 n1986_not ; n1987
g1939 nor n1985 n1987 ; n1988
g1940 and n1984_not n1988 ; n1989
g1941 and n1983_not n1989 ; n1990
g1942 and n1983 n1989_not ; n1991
g1943 nor n1990 n1991 ; n1992
g1944 and n1976_not n1992 ; n1993
g1945 and n1976 n1992_not ; n1994
g1946 and n1013_not n1550 ; n1995
g1947 and n1013 n1549 ; n1996
g1948 and n1130_not n1183 ; n1997
g1949 and n1487 n1997_not ; n1998
g1950 nor n1996 n1998 ; n1999
g1951 and n1995_not n1999 ; n2000
g1952 and n275_not n1368 ; n2001
g1953 and n275 n1317 ; n2002
g1954 and n279 n1371 ; n2003
g1955 and n279_not n1315 ; n2004
g1956 nor n2003 n2004 ; n2005
g1957 and n2002_not n2005 ; n2006
g1958 and n2001_not n2006 ; n2007
g1959 and n2000 n2007_not ; n2008
g1960 and n2000_not n2007 ; n2009
g1961 nor n2008 n2009 ; n2010
g1962 and n1183_not n1550 ; n2011
g1963 and n1183 n1549 ; n2012
g1964 and n275 n1130_not ; n2013
g1965 and n1487 n2013_not ; n2014
g1966 nor n2012 n2014 ; n2015
g1967 and n2011_not n2015 ; n2016
g1968 and n286_not n1368 ; n2017
g1969 and n286 n1177_not ; n2018
g1970 nor n1371 n2018 ; n2019
g1971 and n2017_not n2019 ; n2020
g1972 and n1177 n2020 ; n2021
g1973 and n2016 n2021 ; n2022
g1974 and n2010 n2022_not ; n2023
g1975 and n2010_not n2022 ; n2024
g1976 and n279_not n1368 ; n2025
g1977 and n279 n1317 ; n2026
g1978 and n286_not n1315 ; n2027
g1979 nor n1177 n2020 ; n2028
g1980 and n275_not n1550 ; n2029
g1981 and n275 n1549 ; n2030
g1982 nor n279 n1487 ; n2031
g1983 and n1130 n1487 ; n2032
g1984 and n279 n2032_not ; n2033
g1985 nor n2031 n2033 ; n2034
g1986 nor n2030 n2034 ; n2035
g1987 and n2029_not n2035 ; n2036
g1988 and n286 n1130_not ; n2037
g1989 and n2031_not n2037 ; n2038
g1990 nor n2036 n2038 ; n2039
g1991 nor n2021 n2039 ; n2040
g1992 and n2028_not n2040 ; n2041
g1993 and n2036 n2038 ; n2042
g1994 nor n2041 n2042 ; n2043
g1995 nor n2016 n2021 ; n2044
g1996 nor n2022 n2044 ; n2045
g1997 and n2043 n2045_not ; n2046
g1998 and n286 n1371 ; n2047
g1999 nor n2046 n2047 ; n2048
g2000 and n2027_not n2048 ; n2049
g2001 and n2026_not n2049 ; n2050
g2002 and n2025_not n2050 ; n2051
g2003 and n2043_not n2045 ; n2052
g2004 nor n2051 n2052 ; n2053
g2005 nor n286 n1194 ; n2054
g2006 and n2053 n2054_not ; n2055
g2007 nor n2024 n2055 ; n2056
g2008 and n2023_not n2056 ; n2057
g2009 and n2053_not n2054 ; n2058
g2010 nor n2057 n2058 ; n2059
g2011 and n1959 n1962_not ; n2060
g2012 and n1960_not n1963 ; n2061
g2013 nor n2060 n2061 ; n2062
g2014 and n2059 n2062 ; n2063
g2015 and n2000 n2007 ; n2064
g2016 nor n2024 n2064 ; n2065
g2017 nor n2063 n2065 ; n2066
g2018 nor n2059 n2062 ; n2067
g2019 nor n2066 n2067 ; n2068
g2020 nor n1963 n1968 ; n2069
g2021 nor n1967 n1968 ; n2070
g2022 nor n2069 n2070 ; n2071
g2023 and n2068 n2071 ; n2072
g2024 nor n1994 n2072 ; n2073
g2025 and n1993_not n2073 ; n2074
g2026 nor n2068 n2071 ; n2075
g2027 nor n2074 n2075 ; n2076
g2028 nor n1969 n2076 ; n2077
g2029 and n1969 n2076 ; n2078
g2030 and n1897 n1915_not ; n2079
g2031 nor n1914 n1915 ; n2080
g2032 nor n2079 n2080 ; n2081
g2033 nor n1868 n1873 ; n2082
g2034 nor n1874 n2082 ; n2083
g2035 and n1983 n1989 ; n2084
g2036 nor n1994 n2084 ; n2085
g2037 and n2083 n2085_not ; n2086
g2038 and n2083_not n2085 ; n2087
g2039 nor n2086 n2087 ; n2088
g2040 and n2081_not n2088 ; n2089
g2041 and n2081 n2088_not ; n2090
g2042 nor n2089 n2090 ; n2091
g2043 and n2078_not n2091 ; n2092
g2044 nor n2077 n2092 ; n2093
g2045 nor n2086 n2089 ; n2094
g2046 nor n2093 n2094 ; n2095
g2047 and n2093 n2094 ; n2096
g2048 and n1922_not n1925 ; n2097
g2049 nor n1926 n2097 ; n2098
g2050 and n2096_not n2098 ; n2099
g2051 nor n2095 n2099 ; n2100
g2052 and n1927 n2100 ; n2101
g2053 nor n1890 n2101 ; n2102
g2054 and n1889_not n2102 ; n2103
g2055 nor n1927 n2100 ; n2104
g2056 nor n2103 n2104 ; n2105
g2057 nor n1884 n1890 ; n2106
g2058 nor n2105 n2106 ; n2107
g2059 and n2105 n2106 ; n2108
g2060 and n1850 n1853 ; n2109
g2061 nor n1854 n2109 ; n2110
g2062 and n2108_not n2110 ; n2111
g2063 nor n2107 n2111 ; n2112
g2064 and n1855 n2112 ; n2113
g2065 and n1793 n1796 ; n2114
g2066 nor n2113 n2114 ; n2115
g2067 and n1797_not n2115 ; n2116
g2068 nor n1855 n2112 ; n2117
g2069 nor n2116 n2117 ; n2118
g2070 and n1799 n1801_not ; n2119
g2071 nor n1802 n2119 ; n2120
g2072 and n2118_not n2120 ; n2121
g2073 nor n1802 n2121 ; n2122
g2074 and n1746 n1748_not ; n2123
g2075 nor n1749 n2123 ; n2124
g2076 and n2122_not n2124 ; n2125
g2077 nor n1749 n2125 ; n2126
g2078 and n1666 n1668_not ; n2127
g2079 nor n1669 n2127 ; n2128
g2080 and n2126_not n2128 ; n2129
g2081 nor n1669 n2129 ; n2130
g2082 and n1623 n1625_not ; n2131
g2083 nor n1626 n2131 ; n2132
g2084 and n2130_not n2132 ; n2133
g2085 nor n1626 n2133 ; n2134
g2086 nor n1548 n2134 ; n2135
g2087 nor n1545 n2135 ; n2136
g2088 and n1424 n1427 ; n2137
g2089 nor n1428 n2137 ; n2138
g2090 and n2136_not n2138 ; n2139
g2091 nor n1428 n2139 ; n2140
g2092 nor n1295 n2140 ; n2141
g2093 nor n1292 n2141 ; n2142
g2094 and n1234 n1236_not ; n2143
g2095 nor n1237 n2143 ; n2144
g2096 and n2142_not n2144 ; n2145
g2097 nor n1237 n2145 ; n2146
g2098 nor n1074 n2146 ; n2147
g2099 nor n1068 n1071 ; n2148
g2100 nor n2147 n2148 ; n2149
g2101 and n895 n897_not ; n2150
g2102 nor n898 n2150 ; n2151
g2103 and n2149_not n2151 ; n2152
g2104 nor n898 n2152 ; n2153
g2105 nor n728 n2153 ; n2154
g2106 nor n722 n725 ; n2155
g2107 nor n2154 n2155 ; n2156
g2108 and n683 n2156_not ; n2157
g2109 and n683_not n2156 ; n2158
g2110 nor n2157 n2158 ; n2159
g2111 and n536 n2159 ; n2160
g2112 nor n536 n2159 ; n2161
g2113 nor n2160 n2161 ; n2162
g2114 nor n393 n2162 ; n2163
g2115 and n393 n2162 ; n2164
g2116 nor n134 n468 ; n2165
g2117 and n219_not n2165 ; n2166
g2118 nor n254 n329 ; n2167
g2119 and n358_not n2167 ; n2168
g2120 and n326_not n2168 ; n2169
g2121 and n342_not n2169 ; n2170
g2122 and n760 n2170 ; n2171
g2123 and n226_not n2171 ; n2172
g2124 and n218_not n2172 ; n2173
g2125 and n167_not n2173 ; n2174
g2126 and n206_not n2174 ; n2175
g2127 and n190_not n2175 ; n2176
g2128 and n589_not n2176 ; n2177
g2129 and n736_not n2177 ; n2178
g2130 and n415_not n626 ; n2179
g2131 and n297_not n2179 ; n2180
g2132 and n356_not n2180 ; n2181
g2133 and n361_not n968 ; n2182
g2134 and n142_not n2182 ; n2183
g2135 and n555 n2183 ; n2184
g2136 and n476 n2184 ; n2185
g2137 and n1091 n2185 ; n2186
g2138 and n2181 n2186 ; n2187
g2139 and n986 n2187 ; n2188
g2140 and n753 n2188 ; n2189
g2141 and n154_not n2189 ; n2190
g2142 and n140_not n792 ; n2191
g2143 and n299_not n2191 ; n2192
g2144 and n458_not n2192 ; n2193
g2145 and n357_not n2193 ; n2194
g2146 and n148_not n2194 ; n2195
g2147 and n553_not n2195 ; n2196
g2148 and n153 n808 ; n2197
g2149 and n397 n2197 ; n2198
g2150 and n773 n2198 ; n2199
g2151 and n2196 n2199 ; n2200
g2152 and n2190 n2200 ; n2201
g2153 and n2178 n2201 ; n2202
g2154 and n2166 n2202 ; n2203
g2155 and n328_not n2203 ; n2204
g2156 and n228_not n2204 ; n2205
g2157 and n177_not n2205 ; n2206
g2158 and n504_not n2206 ; n2207
g2159 and n367_not n2207 ; n2208
g2160 and n215_not n2208 ; n2209
g2161 and n728 n2153 ; n2210
g2162 nor n2154 n2210 ; n2211
g2163 nor n2209 n2211 ; n2212
g2164 and n145 n794 ; n2213
g2165 and n319 n2213 ; n2214
g2166 and n474 n2214 ; n2215
g2167 and n637 n2215 ; n2216
g2168 and n739 n2216 ; n2217
g2169 and n967 n2217 ; n2218
g2170 and n606 n2218 ; n2219
g2171 and n1104 n2219 ; n2220
g2172 and n458_not n2220 ; n2221
g2173 and n297_not n2221 ; n2222
g2174 and n358_not n2222 ; n2223
g2175 and n168_not n2223 ; n2224
g2176 and n237_not n2224 ; n2225
g2177 and n2149 n2151_not ; n2226
g2178 nor n2152 n2226 ; n2227
g2179 nor n2225 n2227 ; n2228
g2180 and n2225 n2227 ; n2229
g2181 and n331 n2183 ; n2230
g2182 and n236 n2230 ; n2231
g2183 and n301 n2231 ; n2232
g2184 and n637 n2232 ; n2233
g2185 and n2166 n2233 ; n2234
g2186 and n355 n2234 ; n2235
g2187 and n221_not n2235 ; n2236
g2188 and n394_not n2236 ; n2237
g2189 and n225_not n2237 ; n2238
g2190 and n206_not n2238 ; n2239
g2191 and n254_not n906 ; n2240
g2192 and n447_not n2240 ; n2241
g2193 and n148_not n2241 ; n2242
g2194 and n111_not n2242 ; n2243
g2195 and n238_not n2243 ; n2244
g2196 and n581 n628 ; n2245
g2197 and n2244 n2245 ; n2246
g2198 and n227_not n2246 ; n2247
g2199 and n417_not n2247 ; n2248
g2200 and n123_not n2248 ; n2249
g2201 and n736_not n2249 ; n2250
g2202 nor n178 n506 ; n2251
g2203 and n471_not n2251 ; n2252
g2204 nor n302 n313 ; n2253
g2205 and n445_not n2253 ; n2254
g2206 and n478 n2254 ; n2255
g2207 and n2252 n2255 ; n2256
g2208 and n156 n2256 ; n2257
g2209 and n577 n2257 ; n2258
g2210 and n644 n2258 ; n2259
g2211 and n2250 n2259 ; n2260
g2212 and n2239 n2260 ; n2261
g2213 and n317_not n2261 ; n2262
g2214 and n336_not n2262 ; n2263
g2215 and n554_not n2263 ; n2264
g2216 and n1074 n2146 ; n2265
g2217 nor n2147 n2265 ; n2266
g2218 nor n2264 n2266 ; n2267
g2219 and n396 n2252 ; n2268
g2220 and n451 n2268 ; n2269
g2221 and n139_not n2269 ; n2270
g2222 and n188_not n2270 ; n2271
g2223 and n129_not n2271 ; n2272
g2224 and n359_not n2272 ; n2273
g2225 and n335_not n2273 ; n2274
g2226 and n367_not n2274 ; n2275
g2227 and n599_not n2275 ; n2276
g2228 nor n447 n552 ; n2277
g2229 and n237_not n2277 ; n2278
g2230 and n152_not n2239 ; n2279
g2231 and n296_not n2279 ; n2280
g2232 and n215_not n2280 ; n2281
g2233 and n1459 n2281 ; n2282
g2234 and n2278 n2282 ; n2283
g2235 and n325 n2283 ; n2284
g2236 and n2196 n2284 ; n2285
g2237 and n2276 n2285 ; n2286
g2238 and n980 n2286 ; n2287
g2239 and n176_not n2287 ; n2288
g2240 and n343_not n2288 ; n2289
g2241 and n167_not n2289 ; n2290
g2242 and n360_not n2290 ; n2291
g2243 and n313_not n2291 ; n2292
g2244 and n2142 n2144_not ; n2293
g2245 nor n2145 n2293 ; n2294
g2246 nor n2292 n2294 ; n2295
g2247 and n2292 n2294 ; n2296
g2248 nor n138 n227 ; n2297
g2249 and n123_not n2297 ; n2298
g2250 and n172_not n2298 ; n2299
g2251 and n234_not n2299 ; n2300
g2252 and n357_not n2300 ; n2301
g2253 and n216_not n2301 ; n2302
g2254 and n168_not n2302 ; n2303
g2255 and n141 n1116 ; n2304
g2256 and n944 n2304 ; n2305
g2257 and n644 n2305 ; n2306
g2258 and n369 n2306 ; n2307
g2259 and n337_not n2307 ; n2308
g2260 and n458_not n2308 ; n2309
g2261 and n447_not n2309 ; n2310
g2262 and n347_not n2310 ; n2311
g2263 and n106_not n923 ; n2312
g2264 and n326_not n2312 ; n2313
g2265 nor n217 n228 ; n2314
g2266 and n146_not n2314 ; n2315
g2267 and n211_not n2315 ; n2316
g2268 and n469_not n2316 ; n2317
g2269 and n2313 n2317 ; n2318
g2270 and n2311 n2318 ; n2319
g2271 and n2303 n2319 ; n2320
g2272 and n328_not n2320 ; n2321
g2273 and n408_not n2321 ; n2322
g2274 and n194_not n2322 ; n2323
g2275 and n219_not n2323 ; n2324
g2276 and n298_not n2324 ; n2325
g2277 and n450 n2325 ; n2326
g2278 and n445_not n2326 ; n2327
g2279 and n1295 n2140 ; n2328
g2280 nor n2141 n2328 ; n2329
g2281 nor n2327 n2329 ; n2330
g2282 and n213_not n508 ; n2331
g2283 and n736_not n2331 ; n2332
g2284 and n345_not n2332 ; n2333
g2285 and n303 n759 ; n2334
g2286 and n931 n2334 ; n2335
g2287 and n169_not n2335 ; n2336
g2288 and n114_not n2336 ; n2337
g2289 and n326_not n2337 ; n2338
g2290 and n469_not n2338 ; n2339
g2291 nor n138 n146 ; n2340
g2292 nor n106 n348 ; n2341
g2293 and n238_not n2341 ; n2342
g2294 and n432 n2342 ; n2343
g2295 and n2340 n2343 ; n2344
g2296 and n1106 n2344 ; n2345
g2297 and n344 n2345 ; n2346
g2298 and n314 n2346 ; n2347
g2299 and n2339 n2347 ; n2348
g2300 and n995 n2348 ; n2349
g2301 and n930 n2349 ; n2350
g2302 and n2333 n2350 ; n2351
g2303 and n152_not n2351 ; n2352
g2304 and n217_not n2352 ; n2353
g2305 and n495_not n2353 ; n2354
g2306 and n2136 n2138_not ; n2355
g2307 nor n2139 n2355 ; n2356
g2308 nor n2354 n2356 ; n2357
g2309 and n2354 n2356 ; n2358
g2310 and n141 n312_not ; n2359
g2311 and n417_not n2359 ; n2360
g2312 and n313_not n2360 ; n2361
g2313 and n224_not n2361 ; n2362
g2314 and n553_not n2362 ; n2363
g2315 and n235_not n2363 ; n2364
g2316 nor n255 n449 ; n2365
g2317 and n554_not n2365 ; n2366
g2318 nor n194 n237 ; n2367
g2319 and n2366 n2367 ; n2368
g2320 and n910 n2368 ; n2369
g2321 and n188_not n2369 ; n2370
g2322 and n327_not n2370 ; n2371
g2323 and n348_not n2371 ; n2372
g2324 and n329_not n2372 ; n2373
g2325 and n191_not n2373 ; n2374
g2326 and n503_not n2374 ; n2375
g2327 and n382 n448 ; n2376
g2328 and n2375 n2376 ; n2377
g2329 and n753 n2377 ; n2378
g2330 and n2364 n2378 ; n2379
g2331 and n196_not n2379 ; n2380
g2332 and n221_not n2380 ; n2381
g2333 and n394_not n2381 ; n2382
g2334 and n167_not n2382 ; n2383
g2335 and n347_not n2383 ; n2384
g2336 and n472_not n2384 ; n2385
g2337 and n1548 n2134 ; n2386
g2338 nor n2135 n2386 ; n2387
g2339 nor n2385 n2387 ; n2388
g2340 and n564 n2254 ; n2389
g2341 and n906 n2389 ; n2390
g2342 and n411 n2390 ; n2391
g2343 and n360_not n2391 ; n2392
g2344 and n114_not n2392 ; n2393
g2345 and n326_not n2393 ; n2394
g2346 and n223_not n2394 ; n2395
g2347 and n416 n473 ; n2396
g2348 and n298_not n2396 ; n2397
g2349 and n118_not n2397 ; n2398
g2350 and n224_not n2398 ; n2399
g2351 and n367_not n2399 ; n2400
g2352 and n590 n2400 ; n2401
g2353 and n2395 n2401 ; n2402
g2354 and n752 n2402 ; n2403
g2355 and n986 n2403 ; n2404
g2356 and n149 n2404 ; n2405
g2357 and n228_not n2405 ; n2406
g2358 and n219_not n2406 ; n2407
g2359 and n226_not n2407 ; n2408
g2360 and n336_not n2408 ; n2409
g2361 and n234_not n2409 ; n2410
g2362 and n258_not n2410 ; n2411
g2363 and n554_not n2411 ; n2412
g2364 and n342_not n2412 ; n2413
g2365 and n296_not n2413 ; n2414
g2366 and n2130 n2132_not ; n2415
g2367 nor n2133 n2415 ; n2416
g2368 nor n2414 n2416 ; n2417
g2369 nor n553 n599 ; n2418
g2370 and n335_not n2418 ; n2419
g2371 and n111_not n2419 ; n2420
g2372 and n477_not n2420 ; n2421
g2373 nor n296 n449 ; n2422
g2374 and n970 n2422 ; n2423
g2375 and n2421 n2423 ; n2424
g2376 and n2278 n2424 ; n2425
g2377 and n373 n2425 ; n2426
g2378 and n2333 n2426 ; n2427
g2379 and n926 n2427 ; n2428
g2380 and n359_not n2428 ; n2429
g2381 and n358_not n2429 ; n2430
g2382 and n472_not n2430 ; n2431
g2383 and n223_not n2431 ; n2432
g2384 nor n351 n504 ; n2433
g2385 and n396 n806 ; n2434
g2386 and n2433 n2434 ; n2435
g2387 and n2400 n2435 ; n2436
g2388 and n325 n2436 ; n2437
g2389 and n323 n2437 ; n2438
g2390 and n983 n2438 ; n2439
g2391 and n2432 n2439 ; n2440
g2392 and n165 n2440 ; n2441
g2393 and n328_not n2441 ; n2442
g2394 and n214_not n2442 ; n2443
g2395 and n257_not n2443 ; n2444
g2396 and n360_not n2444 ; n2445
g2397 and n238_not n2445 ; n2446
g2398 and n2126 n2128_not ; n2447
g2399 nor n2129 n2447 ; n2448
g2400 nor n2446 n2448 ; n2449
g2401 and n2446 n2448 ; n2450
g2402 and n152_not n1117 ; n2451
g2403 and n227_not n2451 ; n2452
g2404 and n347_not n2452 ; n2453
g2405 and n554_not n2453 ; n2454
g2406 nor n176 n312 ; n2455
g2407 and n370_not n2455 ; n2456
g2408 and n361_not n2456 ; n2457
g2409 and n132_not n2457 ; n2458
g2410 and n2454 n2458 ; n2459
g2411 and n343_not n2459 ; n2460
g2412 and n458_not n2460 ; n2461
g2413 and n359_not n2461 ; n2462
g2414 and n552_not n2462 ; n2463
g2415 and n154_not n2463 ; n2464
g2416 and n256 n2422 ; n2465
g2417 and n474 n2465 ; n2466
g2418 and n2339 n2466 ; n2467
g2419 and n2464 n2467 ; n2468
g2420 and n789 n2468 ; n2469
g2421 and n337_not n2469 ; n2470
g2422 and n208_not n2470 ; n2471
g2423 and n134_not n2471 ; n2472
g2424 and n192_not n2472 ; n2473
g2425 and n123_not n2473 ; n2474
g2426 and n224_not n2474 ; n2475
g2427 and n357_not n2475 ; n2476
g2428 and n445_not n2476 ; n2477
g2429 and n2122 n2124_not ; n2478
g2430 nor n2125 n2478 ; n2479
g2431 nor n2477 n2479 ; n2480
g2432 and n2477 n2479 ; n2481
g2433 nor n2118 n2121 ; n2482
g2434 and n2120 n2121_not ; n2483
g2435 nor n2482 n2483 ; n2484
g2436 and n777 n1096 ; n2485
g2437 and n914 n2485 ; n2486
g2438 and n373 n2486 ; n2487
g2439 and n2395 n2487 ; n2488
g2440 and n739 n2488 ; n2489
g2441 and n2190 n2489 ; n2490
g2442 and n417_not n2490 ; n2491
g2443 and n192_not n2491 ; n2492
g2444 and n358_not n2492 ; n2493
g2445 and n190_not n2493 ; n2494
g2446 and n599_not n2494 ; n2495
g2447 and n2484_not n2495 ; n2496
g2448 nor n2480 n2496 ; n2497
g2449 and n2481_not n2497 ; n2498
g2450 nor n2480 n2498 ; n2499
g2451 nor n2449 n2499 ; n2500
g2452 and n2450_not n2500 ; n2501
g2453 nor n2449 n2501 ; n2502
g2454 and n2414 n2416 ; n2503
g2455 nor n2417 n2503 ; n2504
g2456 and n2502_not n2504 ; n2505
g2457 nor n2417 n2505 ; n2506
g2458 and n2385 n2387 ; n2507
g2459 nor n2388 n2507 ; n2508
g2460 and n2506_not n2508 ; n2509
g2461 nor n2388 n2509 ; n2510
g2462 nor n2357 n2510 ; n2511
g2463 and n2358_not n2511 ; n2512
g2464 nor n2357 n2512 ; n2513
g2465 nor n2327 n2330 ; n2514
g2466 nor n2329 n2330 ; n2515
g2467 nor n2514 n2515 ; n2516
g2468 nor n2513 n2516 ; n2517
g2469 nor n2330 n2517 ; n2518
g2470 nor n2295 n2518 ; n2519
g2471 and n2296_not n2519 ; n2520
g2472 nor n2295 n2520 ; n2521
g2473 and n2264 n2266 ; n2522
g2474 nor n2267 n2522 ; n2523
g2475 and n2521_not n2523 ; n2524
g2476 nor n2267 n2524 ; n2525
g2477 nor n2228 n2525 ; n2526
g2478 and n2229_not n2526 ; n2527
g2479 nor n2228 n2527 ; n2528
g2480 and n2209 n2211 ; n2529
g2481 nor n2212 n2529 ; n2530
g2482 and n2528_not n2530 ; n2531
g2483 nor n2212 n2531 ; n2532
g2484 nor n2163 n2532 ; n2533
g2485 and n2164_not n2533 ; n2534
g2486 nor n2163 n2534 ; n2535
g2487 and n408_not n796 ; n2536
g2488 and n188_not n2536 ; n2537
g2489 and n227_not n2537 ; n2538
g2490 and n174_not n2538 ; n2539
g2491 and n368_not n2539 ; n2540
g2492 and n478 n1091 ; n2541
g2493 and n2339 n2541 ; n2542
g2494 and n1468 n2542 ; n2543
g2495 and n2540 n2543 ; n2544
g2496 and n653 n2544 ; n2545
g2497 and n149 n2545 ; n2546
g2498 and n299_not n2546 ; n2547
g2499 and n945 n2547 ; n2548
g2500 and n552_not n2548 ; n2549
g2501 and n554_not n2549 ; n2550
g2502 and n223_not n2550 ; n2551
g2503 and n2535 n2551 ; n2552
g2504 nor n2535 n2551 ; n2553
g2505 nor n2552 n2553 ; n2554
g2506 and n295 n2554_not ; n2555
g2507 and n279_not n286 ; n2556
g2508 and n279 n286_not ; n2557
g2509 nor n2556 n2557 ; n2558
g2510 and n282_not n294 ; n2559
g2511 and n2558 n2559 ; n2560
g2512 and n2528 n2530_not ; n2561
g2513 nor n2531 n2561 ; n2562
g2514 and n2560 n2562 ; n2563
g2515 nor n2532 n2534 ; n2564
g2516 and n2164_not n2535 ; n2565
g2517 nor n2564 n2565 ; n2566
g2518 and n294 n2558_not ; n2567
g2519 and n2566_not n2567 ; n2568
g2520 nor n2563 n2568 ; n2569
g2521 and n2555_not n2569 ; n2570
g2522 nor n282 n294 ; n2571
g2523 and n2562 n2566_not ; n2572
g2524 nor n2525 n2527 ; n2573
g2525 and n2229_not n2528 ; n2574
g2526 nor n2573 n2574 ; n2575
g2527 and n2562 n2575_not ; n2576
g2528 and n2521 n2523_not ; n2577
g2529 nor n2524 n2577 ; n2578
g2530 and n2575_not n2578 ; n2579
g2531 nor n2518 n2520 ; n2580
g2532 and n2296_not n2521 ; n2581
g2533 nor n2580 n2581 ; n2582
g2534 and n2578 n2582_not ; n2583
g2535 nor n2513 n2517 ; n2584
g2536 nor n2516 n2517 ; n2585
g2537 nor n2584 n2585 ; n2586
g2538 nor n2582 n2586 ; n2587
g2539 nor n2510 n2512 ; n2588
g2540 and n2358_not n2513 ; n2589
g2541 nor n2588 n2589 ; n2590
g2542 nor n2586 n2590 ; n2591
g2543 and n2506 n2508_not ; n2592
g2544 nor n2509 n2592 ; n2593
g2545 and n2590_not n2593 ; n2594
g2546 and n2502 n2504_not ; n2595
g2547 nor n2505 n2595 ; n2596
g2548 and n2593 n2596 ; n2597
g2549 nor n2499 n2501 ; n2598
g2550 and n2450_not n2502 ; n2599
g2551 nor n2598 n2599 ; n2600
g2552 and n2596 n2600_not ; n2601
g2553 nor n2496 n2498 ; n2602
g2554 and n2481_not n2499 ; n2603
g2555 nor n2602 n2603 ; n2604
g2556 nor n2600 n2604 ; n2605
g2557 and n2484 n2495_not ; n2606
g2558 nor n2496 n2606 ; n2607
g2559 nor n2604 n2607 ; n2608
g2560 and n2600 n2608 ; n2609
g2561 nor n2605 n2609 ; n2610
g2562 and n2596_not n2600 ; n2611
g2563 nor n2610 n2611 ; n2612
g2564 and n2601_not n2612 ; n2613
g2565 nor n2601 n2613 ; n2614
g2566 nor n2593 n2596 ; n2615
g2567 nor n2614 n2615 ; n2616
g2568 and n2597_not n2616 ; n2617
g2569 nor n2597 n2617 ; n2618
g2570 and n2590 n2593_not ; n2619
g2571 nor n2594 n2619 ; n2620
g2572 and n2618_not n2620 ; n2621
g2573 nor n2594 n2621 ; n2622
g2574 and n2586 n2590 ; n2623
g2575 nor n2591 n2623 ; n2624
g2576 and n2622_not n2624 ; n2625
g2577 nor n2591 n2625 ; n2626
g2578 and n2582 n2586 ; n2627
g2579 nor n2587 n2627 ; n2628
g2580 and n2626_not n2628 ; n2629
g2581 nor n2587 n2629 ; n2630
g2582 and n2578_not n2582 ; n2631
g2583 nor n2583 n2631 ; n2632
g2584 and n2630_not n2632 ; n2633
g2585 nor n2583 n2633 ; n2634
g2586 and n2575 n2578_not ; n2635
g2587 nor n2579 n2635 ; n2636
g2588 and n2634_not n2636 ; n2637
g2589 nor n2579 n2637 ; n2638
g2590 and n2562_not n2575 ; n2639
g2591 nor n2576 n2639 ; n2640
g2592 and n2638_not n2640 ; n2641
g2593 nor n2576 n2641 ; n2642
g2594 and n2562_not n2566 ; n2643
g2595 nor n2572 n2643 ; n2644
g2596 and n2642_not n2644 ; n2645
g2597 nor n2572 n2645 ; n2646
g2598 nor n2554 n2566 ; n2647
g2599 and n2554 n2566 ; n2648
g2600 nor n2647 n2648 ; n2649
g2601 and n2646_not n2649 ; n2650
g2602 and n2646 n2649_not ; n2651
g2603 nor n2650 n2651 ; n2652
g2604 and n2571 n2652 ; n2653
g2605 and n2570 n2653_not ; n2654
g2606 nor n275 n2654 ; n2655
g2607 and n275 n2654 ; n2656
g2608 nor n2655 n2656 ; n2657
g2609 and n669 n677_not ; n2658
g2610 and n669_not n677 ; n2659
g2611 nor n2658 n2659 ; n2660
g2612 nor n2607 n2660 ; n2661
g2613 nor n525 n2661 ; n2662
g2614 and n529 n677_not ; n2663
g2615 and n529_not n677 ; n2664
g2616 nor n2663 n2664 ; n2665
g2617 and n2660 n2665_not ; n2666
g2618 and n2607_not n2666 ; n2667
g2619 and n532 n2660_not ; n2668
g2620 and n2604_not n2668 ; n2669
g2621 nor n2667 n2669 ; n2670
g2622 and n2604 n2607_not ; n2671
g2623 and n2604_not n2607 ; n2672
g2624 nor n2671 n2672 ; n2673
g2625 nor n532 n2660 ; n2674
g2626 and n2673_not n2674 ; n2675
g2627 and n2670 n2675_not ; n2676
g2628 nor n525 n2676 ; n2677
g2629 nor n525 n2677 ; n2678
g2630 nor n2676 n2677 ; n2679
g2631 nor n2678 n2679 ; n2680
g2632 and n2662 n2680_not ; n2681
g2633 and n2662_not n2680 ; n2682
g2634 nor n2681 n2682 ; n2683
g2635 and n832 n1021_not ; n2684
g2636 and n832_not n1021 ; n2685
g2637 nor n2684 n2685 ; n2686
g2638 and n669 n840_not ; n2687
g2639 and n669_not n840 ; n2688
g2640 nor n2687 n2688 ; n2689
g2641 nor n2686 n2689 ; n2690
g2642 and n832 n840_not ; n2691
g2643 and n832_not n840 ; n2692
g2644 nor n2691 n2692 ; n2693
g2645 and n2686 n2689_not ; n2694
g2646 and n2693 n2694 ; n2695
g2647 and n2600_not n2695 ; n2696
g2648 and n2686 n2693_not ; n2697
g2649 and n2596 n2697 ; n2698
g2650 and n2686_not n2689 ; n2699
g2651 and n2593 n2699 ; n2700
g2652 nor n2698 n2700 ; n2701
g2653 and n2696_not n2701 ; n2702
g2654 and n2690_not n2702 ; n2703
g2655 nor n2614 n2617 ; n2704
g2656 and n2615_not n2618 ; n2705
g2657 nor n2704 n2705 ; n2706
g2658 and n2702 n2706 ; n2707
g2659 nor n2703 n2707 ; n2708
g2660 and n669 n2708_not ; n2709
g2661 and n669_not n2708 ; n2710
g2662 nor n2709 n2710 ; n2711
g2663 and n2683 n2711 ; n2712
g2664 nor n2607 n2686 ; n2713
g2665 nor n669 n2713 ; n2714
g2666 and n2607_not n2697 ; n2715
g2667 and n2604_not n2699 ; n2716
g2668 nor n2715 n2716 ; n2717
g2669 and n2673_not n2690 ; n2718
g2670 and n2717 n2718_not ; n2719
g2671 nor n669 n2719 ; n2720
g2672 and n669 n2719 ; n2721
g2673 nor n2720 n2721 ; n2722
g2674 and n2714 n2722 ; n2723
g2675 and n2600_not n2699 ; n2724
g2676 and n2607_not n2695 ; n2725
g2677 and n2604_not n2697 ; n2726
g2678 nor n2725 n2726 ; n2727
g2679 and n2724_not n2727 ; n2728
g2680 and n2690_not n2728 ; n2729
g2681 and n2600 n2672_not ; n2730
g2682 and n2600_not n2672 ; n2731
g2683 nor n2730 n2731 ; n2732
g2684 and n2728 n2732_not ; n2733
g2685 nor n2729 n2733 ; n2734
g2686 and n669 n2734_not ; n2735
g2687 and n669_not n2734 ; n2736
g2688 nor n2735 n2736 ; n2737
g2689 and n2723 n2737 ; n2738
g2690 and n2661 n2738 ; n2739
g2691 and n2738 n2739_not ; n2740
g2692 and n2661 n2739_not ; n2741
g2693 nor n2740 n2741 ; n2742
g2694 and n2600_not n2697 ; n2743
g2695 and n2596 n2699 ; n2744
g2696 and n2604_not n2695 ; n2745
g2697 nor n2744 n2745 ; n2746
g2698 and n2743_not n2746 ; n2747
g2699 nor n2610 n2613 ; n2748
g2700 and n2611_not n2614 ; n2749
g2701 nor n2748 n2749 ; n2750
g2702 and n2690 n2750_not ; n2751
g2703 and n2747 n2751_not ; n2752
g2704 nor n669 n2752 ; n2753
g2705 and n669 n2752 ; n2754
g2706 nor n2753 n2754 ; n2755
g2707 and n2742_not n2755 ; n2756
g2708 nor n2739 n2756 ; n2757
g2709 nor n2683 n2711 ; n2758
g2710 nor n2712 n2758 ; n2759
g2711 and n2757_not n2759 ; n2760
g2712 nor n2712 n2760 ; n2761
g2713 and n2590_not n2699 ; n2762
g2714 and n2596 n2695 ; n2763
g2715 and n2593 n2697 ; n2764
g2716 nor n2763 n2764 ; n2765
g2717 and n2762_not n2765 ; n2766
g2718 and n2618 n2620_not ; n2767
g2719 nor n2621 n2767 ; n2768
g2720 and n2690 n2768 ; n2769
g2721 and n2766 n2769_not ; n2770
g2722 nor n669 n2770 ; n2771
g2723 and n669 n2770 ; n2772
g2724 nor n2771 n2772 ; n2773
g2725 and n2600_not n2668 ; n2774
g2726 and n532_not n2660 ; n2775
g2727 and n2665 n2775 ; n2776
g2728 and n2607_not n2776 ; n2777
g2729 and n2604_not n2666 ; n2778
g2730 nor n2777 n2778 ; n2779
g2731 and n2774_not n2779 ; n2780
g2732 and n2674_not n2780 ; n2781
g2733 and n2732_not n2780 ; n2782
g2734 nor n2781 n2782 ; n2783
g2735 and n525 n2783_not ; n2784
g2736 and n525_not n2783 ; n2785
g2737 nor n2784 n2785 ; n2786
g2738 and n2681 n2786 ; n2787
g2739 nor n2681 n2786 ; n2788
g2740 nor n2787 n2788 ; n2789
g2741 and n2773 n2789 ; n2790
g2742 nor n2773 n2789 ; n2791
g2743 nor n2790 n2791 ; n2792
g2744 and n2761 n2792_not ; n2793
g2745 and n2761_not n2792 ; n2794
g2746 nor n2793 n2794 ; n2795
g2747 and n1013 n1021_not ; n2796
g2748 and n1013_not n1021 ; n2797
g2749 nor n2796 n2797 ; n2798
g2750 and n275 n1183_not ; n2799
g2751 and n275_not n1183 ; n2800
g2752 nor n2799 n2800 ; n2801
g2753 and n2798 n2801_not ; n2802
g2754 and n2578 n2802 ; n2803
g2755 and n1013 n1183_not ; n2804
g2756 and n1013_not n1183 ; n2805
g2757 nor n2804 n2805 ; n2806
g2758 and n2798_not n2801 ; n2807
g2759 and n2806 n2807 ; n2808
g2760 and n2586_not n2808 ; n2809
g2761 and n2801 n2806_not ; n2810
g2762 and n2582_not n2810 ; n2811
g2763 nor n2809 n2811 ; n2812
g2764 and n2803_not n2812 ; n2813
g2765 and n2630 n2632_not ; n2814
g2766 nor n2633 n2814 ; n2815
g2767 and n2813 n2815_not ; n2816
g2768 nor n2798 n2801 ; n2817
g2769 and n2813 n2817_not ; n2818
g2770 nor n2816 n2818 ; n2819
g2771 and n1021 n2819_not ; n2820
g2772 and n1021_not n2819 ; n2821
g2773 nor n2820 n2821 ; n2822
g2774 and n2795 n2822 ; n2823
g2775 and n2582_not n2802 ; n2824
g2776 and n2590_not n2808 ; n2825
g2777 and n2586_not n2810 ; n2826
g2778 nor n2825 n2826 ; n2827
g2779 and n2824_not n2827 ; n2828
g2780 and n2626 n2628_not ; n2829
g2781 nor n2629 n2829 ; n2830
g2782 and n2817 n2830 ; n2831
g2783 and n2828 n2831_not ; n2832
g2784 nor n1021 n2832 ; n2833
g2785 nor n2832 n2833 ; n2834
g2786 nor n1021 n2833 ; n2835
g2787 nor n2834 n2835 ; n2836
g2788 and n2757 n2759_not ; n2837
g2789 nor n2760 n2837 ; n2838
g2790 and n2836_not n2838 ; n2839
g2791 nor n2742 n2756 ; n2840
g2792 and n2755 n2756_not ; n2841
g2793 nor n2840 n2841 ; n2842
g2794 and n2586_not n2802 ; n2843
g2795 and n2593 n2808 ; n2844
g2796 and n2590_not n2810 ; n2845
g2797 nor n2844 n2845 ; n2846
g2798 and n2843_not n2846 ; n2847
g2799 and n2622 n2624_not ; n2848
g2800 nor n2625 n2848 ; n2849
g2801 and n2847 n2849_not ; n2850
g2802 and n2817_not n2847 ; n2851
g2803 nor n2850 n2851 ; n2852
g2804 and n1021 n2852_not ; n2853
g2805 and n1021_not n2852 ; n2854
g2806 nor n2853 n2854 ; n2855
g2807 and n2842_not n2855 ; n2856
g2808 and n2590_not n2802 ; n2857
g2809 and n2596 n2808 ; n2858
g2810 and n2593 n2810 ; n2859
g2811 nor n2858 n2859 ; n2860
g2812 and n2857_not n2860 ; n2861
g2813 and n2768 n2817 ; n2862
g2814 and n2861 n2862_not ; n2863
g2815 nor n1021 n2863 ; n2864
g2816 nor n2863 n2864 ; n2865
g2817 nor n1021 n2864 ; n2866
g2818 nor n2865 n2866 ; n2867
g2819 nor n2723 n2737 ; n2868
g2820 nor n2738 n2868 ; n2869
g2821 and n2867_not n2869 ; n2870
g2822 nor n2714 n2722 ; n2871
g2823 nor n2723 n2871 ; n2872
g2824 and n2600_not n2808 ; n2873
g2825 and n2596 n2810 ; n2874
g2826 and n2593 n2802 ; n2875
g2827 nor n2874 n2875 ; n2876
g2828 and n2873_not n2876 ; n2877
g2829 and n2817_not n2877 ; n2878
g2830 and n2706 n2877 ; n2879
g2831 nor n2878 n2879 ; n2880
g2832 and n1021 n2880_not ; n2881
g2833 and n1021_not n2880 ; n2882
g2834 nor n2881 n2882 ; n2883
g2835 and n2872 n2883 ; n2884
g2836 and n2607_not n2810 ; n2885
g2837 and n2604_not n2802 ; n2886
g2838 nor n2885 n2886 ; n2887
g2839 and n2673_not n2817 ; n2888
g2840 and n2887 n2888_not ; n2889
g2841 nor n1021 n2889 ; n2890
g2842 nor n1021 n2890 ; n2891
g2843 nor n2889 n2890 ; n2892
g2844 nor n2891 n2892 ; n2893
g2845 nor n2607 n2801 ; n2894
g2846 nor n1021 n2894 ; n2895
g2847 and n2893_not n2895 ; n2896
g2848 and n2600_not n2802 ; n2897
g2849 and n2607_not n2808 ; n2898
g2850 and n2604_not n2810 ; n2899
g2851 nor n2898 n2899 ; n2900
g2852 and n2897_not n2900 ; n2901
g2853 and n2732_not n2901 ; n2902
g2854 and n2817_not n2901 ; n2903
g2855 nor n2902 n2903 ; n2904
g2856 and n1021 n2904_not ; n2905
g2857 and n1021_not n2904 ; n2906
g2858 nor n2905 n2906 ; n2907
g2859 and n2896 n2907 ; n2908
g2860 and n2713 n2908 ; n2909
g2861 and n2908 n2909_not ; n2910
g2862 and n2713 n2909_not ; n2911
g2863 nor n2910 n2911 ; n2912
g2864 and n2600_not n2810 ; n2913
g2865 and n2596 n2802 ; n2914
g2866 and n2604_not n2808 ; n2915
g2867 nor n2914 n2915 ; n2916
g2868 and n2913_not n2916 ; n2917
g2869 and n2750_not n2817 ; n2918
g2870 and n2917 n2918_not ; n2919
g2871 nor n1021 n2919 ; n2920
g2872 nor n1021 n2920 ; n2921
g2873 nor n2919 n2920 ; n2922
g2874 nor n2921 n2922 ; n2923
g2875 nor n2912 n2923 ; n2924
g2876 nor n2909 n2924 ; n2925
g2877 nor n2872 n2883 ; n2926
g2878 nor n2884 n2926 ; n2927
g2879 and n2925_not n2927 ; n2928
g2880 nor n2884 n2928 ; n2929
g2881 nor n2867 n2870 ; n2930
g2882 and n2869 n2870_not ; n2931
g2883 nor n2930 n2931 ; n2932
g2884 nor n2929 n2932 ; n2933
g2885 nor n2870 n2933 ; n2934
g2886 nor n2842 n2856 ; n2935
g2887 and n2855 n2856_not ; n2936
g2888 nor n2935 n2936 ; n2937
g2889 nor n2934 n2937 ; n2938
g2890 nor n2856 n2938 ; n2939
g2891 nor n2836 n2839 ; n2940
g2892 and n2838 n2839_not ; n2941
g2893 nor n2940 n2941 ; n2942
g2894 nor n2939 n2942 ; n2943
g2895 nor n2839 n2943 ; n2944
g2896 and n2795 n2823_not ; n2945
g2897 and n2822 n2823_not ; n2946
g2898 nor n2945 n2946 ; n2947
g2899 nor n2944 n2947 ; n2948
g2900 nor n2823 n2948 ; n2949
g2901 and n2586_not n2699 ; n2950
g2902 and n2593 n2695 ; n2951
g2903 and n2590_not n2697 ; n2952
g2904 nor n2951 n2952 ; n2953
g2905 and n2950_not n2953 ; n2954
g2906 and n2690 n2849 ; n2955
g2907 and n2954 n2955_not ; n2956
g2908 nor n669 n2956 ; n2957
g2909 and n669 n2956 ; n2958
g2910 nor n2957 n2958 ; n2959
g2911 and n2600_not n2666 ; n2960
g2912 and n2596 n2668 ; n2961
g2913 and n2604_not n2776 ; n2962
g2914 nor n2961 n2962 ; n2963
g2915 and n2960_not n2963 ; n2964
g2916 and n2674 n2750_not ; n2965
g2917 and n2964 n2965_not ; n2966
g2918 nor n525 n2966 ; n2967
g2919 nor n2966 n2967 ; n2968
g2920 nor n525 n2967 ; n2969
g2921 nor n2968 n2969 ; n2970
g2922 nor n525 n2607 ; n2971
g2923 nor n2787 n2971 ; n2972
g2924 and n2787 n2971 ; n2973
g2925 nor n2970 n2973 ; n2974
g2926 and n2972_not n2974 ; n2975
g2927 nor n2970 n2975 ; n2976
g2928 nor n2973 n2975 ; n2977
g2929 and n2972_not n2977 ; n2978
g2930 nor n2976 n2978 ; n2979
g2931 and n2959 n2979_not ; n2980
g2932 and n2959 n2980_not ; n2981
g2933 nor n2979 n2980 ; n2982
g2934 nor n2981 n2982 ; n2983
g2935 nor n2790 n2794 ; n2984
g2936 and n2983 n2984 ; n2985
g2937 nor n2983 n2984 ; n2986
g2938 nor n2985 n2986 ; n2987
g2939 and n2634 n2636_not ; n2988
g2940 nor n2637 n2988 ; n2989
g2941 and n2575_not n2802 ; n2990
g2942 and n2582_not n2808 ; n2991
g2943 and n2578 n2810 ; n2992
g2944 nor n2991 n2992 ; n2993
g2945 and n2990_not n2993 ; n2994
g2946 and n2989_not n2994 ; n2995
g2947 and n2817_not n2994 ; n2996
g2948 nor n2995 n2996 ; n2997
g2949 and n1021 n2997_not ; n2998
g2950 and n1021_not n2997 ; n2999
g2951 nor n2998 n2999 ; n3000
g2952 and n2987 n3000 ; n3001
g2953 and n2987 n3001_not ; n3002
g2954 and n3000 n3001_not ; n3003
g2955 nor n3002 n3003 ; n3004
g2956 nor n2949 n3004 ; n3005
g2957 nor n2949 n3005 ; n3006
g2958 nor n3004 n3005 ; n3007
g2959 nor n3006 n3007 ; n3008
g2960 and n2657 n3008_not ; n3009
g2961 and n2657 n3009_not ; n3010
g2962 nor n3008 n3009 ; n3011
g2963 nor n3010 n3011 ; n3012
g2964 nor n2944 n2948 ; n3013
g2965 nor n2947 n2948 ; n3014
g2966 nor n3013 n3014 ; n3015
g2967 and n295 n2566_not ; n3016
g2968 and n2560 n2575_not ; n3017
g2969 and n2562 n2567 ; n3018
g2970 nor n3017 n3018 ; n3019
g2971 and n3016_not n3019 ; n3020
g2972 and n2642 n2644_not ; n3021
g2973 nor n2645 n3021 ; n3022
g2974 and n2571 n3022 ; n3023
g2975 and n3020 n3023_not ; n3024
g2976 nor n275 n3024 ; n3025
g2977 and n275 n3024 ; n3026
g2978 nor n3025 n3026 ; n3027
g2979 and n3015_not n3027 ; n3028
g2980 and n3027 n3028_not ; n3029
g2981 nor n3015 n3028 ; n3030
g2982 nor n3029 n3030 ; n3031
g2983 and n2939_not n2942 ; n3032
g2984 and n2939 n2942_not ; n3033
g2985 nor n3032 n3033 ; n3034
g2986 and n295 n2562 ; n3035
g2987 and n2560 n2578 ; n3036
g2988 and n2567 n2575_not ; n3037
g2989 nor n3036 n3037 ; n3038
g2990 and n3035_not n3038 ; n3039
g2991 and n2571_not n3039 ; n3040
g2992 and n2638 n2640_not ; n3041
g2993 nor n2641 n3041 ; n3042
g2994 and n3039 n3042_not ; n3043
g2995 nor n3040 n3043 ; n3044
g2996 and n275 n3044_not ; n3045
g2997 and n275_not n3044 ; n3046
g2998 nor n3045 n3046 ; n3047
g2999 and n3034_not n3047 ; n3048
g3000 nor n2934 n2938 ; n3049
g3001 nor n2937 n2938 ; n3050
g3002 nor n3049 n3050 ; n3051
g3003 and n295 n2575_not ; n3052
g3004 and n2560 n2582_not ; n3053
g3005 and n2567 n2578 ; n3054
g3006 nor n3053 n3054 ; n3055
g3007 and n3052_not n3055 ; n3056
g3008 and n2571_not n3056 ; n3057
g3009 and n2989_not n3056 ; n3058
g3010 nor n3057 n3058 ; n3059
g3011 and n275 n3059_not ; n3060
g3012 and n275_not n3059 ; n3061
g3013 nor n3060 n3061 ; n3062
g3014 and n3051_not n3062 ; n3063
g3015 and n2929_not n2932 ; n3064
g3016 and n2929 n2932_not ; n3065
g3017 nor n3064 n3065 ; n3066
g3018 and n295 n2578 ; n3067
g3019 and n2560 n2586_not ; n3068
g3020 and n2567 n2582_not ; n3069
g3021 nor n3068 n3069 ; n3070
g3022 and n3067_not n3070 ; n3071
g3023 and n2571_not n3071 ; n3072
g3024 and n2815_not n3071 ; n3073
g3025 nor n3072 n3073 ; n3074
g3026 and n275 n3074_not ; n3075
g3027 and n275_not n3074 ; n3076
g3028 nor n3075 n3076 ; n3077
g3029 and n3066_not n3077 ; n3078
g3030 and n295 n2582_not ; n3079
g3031 and n2560 n2590_not ; n3080
g3032 and n2567 n2586_not ; n3081
g3033 nor n3080 n3081 ; n3082
g3034 and n3079_not n3082 ; n3083
g3035 and n2571 n2830 ; n3084
g3036 and n3083 n3084_not ; n3085
g3037 nor n275 n3085 ; n3086
g3038 and n275 n3085 ; n3087
g3039 nor n3086 n3087 ; n3088
g3040 and n2925 n2927_not ; n3089
g3041 nor n2928 n3089 ; n3090
g3042 and n3088 n3090 ; n3091
g3043 nor n2912 n2924 ; n3092
g3044 nor n2923 n2924 ; n3093
g3045 nor n3092 n3093 ; n3094
g3046 and n295 n2586_not ; n3095
g3047 and n2560 n2593 ; n3096
g3048 and n2567 n2590_not ; n3097
g3049 nor n3096 n3097 ; n3098
g3050 and n3095_not n3098 ; n3099
g3051 and n2571_not n3099 ; n3100
g3052 and n2849_not n3099 ; n3101
g3053 nor n3100 n3101 ; n3102
g3054 and n275 n3102_not ; n3103
g3055 and n275_not n3102 ; n3104
g3056 nor n3103 n3104 ; n3105
g3057 and n3094_not n3105 ; n3106
g3058 and n295 n2590_not ; n3107
g3059 and n2560 n2596 ; n3108
g3060 and n2567 n2593 ; n3109
g3061 nor n3108 n3109 ; n3110
g3062 and n3107_not n3110 ; n3111
g3063 and n2571 n2768 ; n3112
g3064 and n3111 n3112_not ; n3113
g3065 nor n275 n3113 ; n3114
g3066 and n275 n3113 ; n3115
g3067 nor n3114 n3115 ; n3116
g3068 nor n2896 n2907 ; n3117
g3069 nor n2908 n3117 ; n3118
g3070 and n3116 n3118 ; n3119
g3071 and n2893 n2895_not ; n3120
g3072 nor n2896 n3120 ; n3121
g3073 and n2560 n2600_not ; n3122
g3074 and n2567 n2596 ; n3123
g3075 and n295 n2593 ; n3124
g3076 nor n3123 n3124 ; n3125
g3077 and n3122_not n3125 ; n3126
g3078 and n2571_not n3126 ; n3127
g3079 and n2706 n3126 ; n3128
g3080 nor n3127 n3128 ; n3129
g3081 and n275 n3129_not ; n3130
g3082 and n275_not n3129 ; n3131
g3083 nor n3130 n3131 ; n3132
g3084 and n3121 n3132 ; n3133
g3085 nor n294 n2607 ; n3134
g3086 nor n275 n3134 ; n3135
g3087 and n2567 n2607_not ; n3136
g3088 and n295 n2604_not ; n3137
g3089 nor n3136 n3137 ; n3138
g3090 and n2571 n2673_not ; n3139
g3091 and n3138 n3139_not ; n3140
g3092 nor n275 n3140 ; n3141
g3093 and n275 n3140 ; n3142
g3094 nor n3141 n3142 ; n3143
g3095 and n3135 n3143 ; n3144
g3096 and n295 n2600_not ; n3145
g3097 and n2560 n2607_not ; n3146
g3098 and n2567 n2604_not ; n3147
g3099 nor n3146 n3147 ; n3148
g3100 and n3145_not n3148 ; n3149
g3101 and n2571_not n3149 ; n3150
g3102 and n2732_not n3149 ; n3151
g3103 nor n3150 n3151 ; n3152
g3104 and n275 n3152_not ; n3153
g3105 and n275_not n3152 ; n3154
g3106 nor n3153 n3154 ; n3155
g3107 and n3144 n3155 ; n3156
g3108 and n2894 n3156 ; n3157
g3109 and n3156 n3157_not ; n3158
g3110 and n2894 n3157_not ; n3159
g3111 nor n3158 n3159 ; n3160
g3112 and n2567 n2600_not ; n3161
g3113 and n295 n2596 ; n3162
g3114 and n2560 n2604_not ; n3163
g3115 nor n3162 n3163 ; n3164
g3116 and n3161_not n3164 ; n3165
g3117 and n2571 n2750_not ; n3166
g3118 and n3165 n3166_not ; n3167
g3119 nor n275 n3167 ; n3168
g3120 and n275 n3167 ; n3169
g3121 nor n3168 n3169 ; n3170
g3122 and n3160_not n3170 ; n3171
g3123 nor n3157 n3171 ; n3172
g3124 nor n3121 n3132 ; n3173
g3125 nor n3133 n3173 ; n3174
g3126 and n3172_not n3174 ; n3175
g3127 nor n3133 n3175 ; n3176
g3128 nor n3116 n3118 ; n3177
g3129 nor n3119 n3177 ; n3178
g3130 and n3176_not n3178 ; n3179
g3131 nor n3119 n3179 ; n3180
g3132 nor n3094 n3106 ; n3181
g3133 and n3105 n3106_not ; n3182
g3134 nor n3181 n3182 ; n3183
g3135 nor n3180 n3183 ; n3184
g3136 nor n3106 n3184 ; n3185
g3137 nor n3088 n3090 ; n3186
g3138 nor n3091 n3186 ; n3187
g3139 and n3185_not n3187 ; n3188
g3140 nor n3091 n3188 ; n3189
g3141 nor n3066 n3078 ; n3190
g3142 and n3077 n3078_not ; n3191
g3143 nor n3190 n3191 ; n3192
g3144 nor n3189 n3192 ; n3193
g3145 nor n3078 n3193 ; n3194
g3146 nor n3051 n3063 ; n3195
g3147 and n3062 n3063_not ; n3196
g3148 nor n3195 n3196 ; n3197
g3149 nor n3194 n3197 ; n3198
g3150 nor n3063 n3198 ; n3199
g3151 and n3034 n3047_not ; n3200
g3152 nor n3048 n3200 ; n3201
g3153 and n3199_not n3201 ; n3202
g3154 nor n3048 n3202 ; n3203
g3155 nor n3031 n3203 ; n3204
g3156 nor n3028 n3204 ; n3205
g3157 and n3012 n3205 ; n3206
g3158 nor n3012 n3205 ; n3207
g3159 nor n3206 n3207 ; n3208
g3160 and a[0] a[22]_not ; n3209
g3161 and a[1] n3209_not ; n3210
g3162 and a[1]_not n3209 ; n3211
g3163 nor n3210 n3211 ; n3212
g3164 and n291_not n3212 ; n3213
g3165 and n291 n3212_not ; n3214
g3166 nor n3213 n3214 ; n3215
g3167 and a[0] n3215_not ; n3216
g3168 and a[0] n3215 ; n3217
g3169 and n324_not n809 ; n3218
g3170 and n485 n3218 ; n3219
g3171 and n431 n3219 ; n3220
g3172 and n2244 n3220 ; n3221
g3173 and n2333 n3221 ; n3222
g3174 and n2418 n3222 ; n3223
g3175 and n976 n3223 ; n3224
g3176 and n504_not n3224 ; n3225
g3177 and n297_not n3225 ; n3226
g3178 and n212_not n3226 ; n3227
g3179 and n258_not n3227 ; n3228
g3180 and n237_not n3228 ; n3229
g3181 and n300_not n808 ; n3230
g3182 and n326_not n3230 ; n3231
g3183 and n200 n3231 ; n3232
g3184 and n2166 n3232 ; n3233
g3185 and n415_not n3233 ; n3234
g3186 and n226_not n3234 ; n3235
g3187 and n213_not n3235 ; n3236
g3188 and n370_not n3236 ; n3237
g3189 and n447_not n3237 ; n3238
g3190 and n335_not n3238 ; n3239
g3191 and n114_not n3239 ; n3240
g3192 and n358_not n3240 ; n3241
g3193 and n106_not n3241 ; n3242
g3194 and n342_not n3242 ; n3243
g3195 and n744 n2366 ; n3244
g3196 and n156 n3244 ; n3245
g3197 and n768 n3245 ; n3246
g3198 and n3243 n3246 ; n3247
g3199 and n210 n3247 ; n3248
g3200 and n150_not n3248 ; n3249
g3201 and n176_not n3249 ; n3250
g3202 and n220_not n3250 ; n3251
g3203 and n227_not n3251 ; n3252
g3204 and n186_not n3252 ; n3253
g3205 and n446_not n3253 ; n3254
g3206 and n361_not n3254 ; n3255
g3207 and n477_not n3255 ; n3256
g3208 and n2552 n3256 ; n3257
g3209 and n3229 n3257 ; n3258
g3210 nor n134 n405 ; n3259
g3211 and n349 n423 ; n3260
g3212 and n1165 n3260 ; n3261
g3213 and n397 n3261 ; n3262
g3214 and n437 n3262 ; n3263
g3215 and n314 n3263 ; n3264
g3216 and n485 n3264 ; n3265
g3217 and n502 n3265 ; n3266
g3218 and n453 n3266 ; n3267
g3219 and n3259 n3267 ; n3268
g3220 and n140_not n3268 ; n3269
g3221 and n3258_not n3269 ; n3270
g3222 and n3258 n3269_not ; n3271
g3223 nor n3270 n3271 ; n3272
g3224 and n3217 n3272 ; n3273
g3225 and n288 n3215_not ; n3274
g3226 and n2552_not n3256 ; n3275
g3227 and n2552 n3256_not ; n3276
g3228 nor n3275 n3276 ; n3277
g3229 and n3274 n3277 ; n3278
g3230 nor n3229 n3257 ; n3279
g3231 nor n3258 n3279 ; n3280
g3232 nor a[0] n3212 ; n3281
g3233 and n3280_not n3281 ; n3282
g3234 nor n3278 n3282 ; n3283
g3235 and n3273_not n3283 ; n3284
g3236 and n3216_not n3284 ; n3285
g3237 and n3277 n3280_not ; n3286
g3238 and n2554_not n3277 ; n3287
g3239 nor n2647 n2650 ; n3288
g3240 and n2554 n3277_not ; n3289
g3241 nor n3287 n3289 ; n3290
g3242 and n3288_not n3290 ; n3291
g3243 nor n3287 n3291 ; n3292
g3244 and n3277_not n3280 ; n3293
g3245 nor n3286 n3293 ; n3294
g3246 and n3292_not n3294 ; n3295
g3247 nor n3286 n3295 ; n3296
g3248 and n3272_not n3280 ; n3297
g3249 and n3272 n3280_not ; n3298
g3250 nor n3297 n3298 ; n3299
g3251 and n3296_not n3299 ; n3300
g3252 and n3296 n3299_not ; n3301
g3253 nor n3300 n3301 ; n3302
g3254 and n3284 n3302_not ; n3303
g3255 nor n3285 n3303 ; n3304
g3256 and n291 n3304_not ; n3305
g3257 and n291_not n3304 ; n3306
g3258 nor n3305 n3306 ; n3307
g3259 and n3208 n3307 ; n3308
g3260 and n3031 n3203 ; n3309
g3261 nor n3204 n3309 ; n3310
g3262 and n3217 n3280_not ; n3311
g3263 and n2554_not n3274 ; n3312
g3264 and n3277 n3281 ; n3313
g3265 nor n3312 n3313 ; n3314
g3266 and n3311_not n3314 ; n3315
g3267 and n3216_not n3315 ; n3316
g3268 and n3292 n3294_not ; n3317
g3269 nor n3295 n3317 ; n3318
g3270 and n3315 n3318_not ; n3319
g3271 nor n3316 n3319 ; n3320
g3272 and n291 n3320_not ; n3321
g3273 and n291_not n3320 ; n3322
g3274 nor n3321 n3322 ; n3323
g3275 and n3310 n3323 ; n3324
g3276 and n3199 n3201_not ; n3325
g3277 and n3217 n3277 ; n3326
g3278 and n2566_not n3274 ; n3327
g3279 and n2554_not n3281 ; n3328
g3280 nor n3327 n3328 ; n3329
g3281 and n3326_not n3329 ; n3330
g3282 and n3288 n3290_not ; n3331
g3283 nor n3291 n3331 ; n3332
g3284 and n3216 n3332 ; n3333
g3285 and n3330 n3333_not ; n3334
g3286 nor n291 n3334 ; n3335
g3287 nor n3334 n3335 ; n3336
g3288 nor n291 n3335 ; n3337
g3289 nor n3336 n3337 ; n3338
g3290 and n2562 n3217 ; n3339
g3291 and n2578 n3274 ; n3340
g3292 and n2575_not n3281 ; n3341
g3293 nor n3340 n3341 ; n3342
g3294 and n3339_not n3342 ; n3343
g3295 nor n291 n3343 ; n3344
g3296 and n3042 n3216 ; n3345
g3297 and n3343 n3345_not ; n3346
g3298 and n291 n3346 ; n3347
g3299 and n291_not n3216 ; n3348
g3300 and n3042 n3348 ; n3349
g3301 and n2575_not n3217 ; n3350
g3302 and n2582_not n3274 ; n3351
g3303 and n2578 n3281 ; n3352
g3304 nor n3351 n3352 ; n3353
g3305 and n3350_not n3353 ; n3354
g3306 nor n291 n3354 ; n3355
g3307 and n2989 n3216 ; n3356
g3308 and n3354 n3356_not ; n3357
g3309 and n291 n3357 ; n3358
g3310 and n2989 n3348 ; n3359
g3311 and n2578 n3217 ; n3360
g3312 and n2586_not n3274 ; n3361
g3313 and n2582_not n3281 ; n3362
g3314 nor n3361 n3362 ; n3363
g3315 and n3360_not n3363 ; n3364
g3316 nor n291 n3364 ; n3365
g3317 and n2815 n3216 ; n3366
g3318 and n3364 n3366_not ; n3367
g3319 and n291 n3367 ; n3368
g3320 and n2815 n3348 ; n3369
g3321 and n3172 n3174_not ; n3370
g3322 and n2586_not n3217 ; n3371
g3323 and n2593 n3274 ; n3372
g3324 and n2590_not n3281 ; n3373
g3325 nor n3372 n3373 ; n3374
g3326 and n3371_not n3374 ; n3375
g3327 nor n291 n3375 ; n3376
g3328 and n2849 n3216 ; n3377
g3329 and n3375 n3377_not ; n3378
g3330 and n291 n3378 ; n3379
g3331 and n2849 n3348 ; n3380
g3332 nor n3144 n3155 ; n3381
g3333 and n2600_not n3274 ; n3382
g3334 and n2596 n3281 ; n3383
g3335 and n2593 n3217 ; n3384
g3336 nor n3383 n3384 ; n3385
g3337 and n3382_not n3385 ; n3386
g3338 nor n291 n3386 ; n3387
g3339 and n2706_not n3216 ; n3388
g3340 and n3386 n3388_not ; n3389
g3341 and n291 n3389 ; n3390
g3342 and n2706_not n3348 ; n3391
g3343 and a[0] n2607_not ; n3392
g3344 and n2732 n3348 ; n3393
g3345 and n2600_not n3217 ; n3394
g3346 and n2607_not n3274 ; n3395
g3347 and n2604_not n3281 ; n3396
g3348 nor n3395 n3396 ; n3397
g3349 and n3394_not n3397 ; n3398
g3350 nor n291 n3398 ; n3399
g3351 and n2673_not n3348 ; n3400
g3352 and n2604_not n3217 ; n3401
g3353 and n2607_not n3281 ; n3402
g3354 nor n291 n3402 ; n3403
g3355 and n3401_not n3403 ; n3404
g3356 and n3400_not n3404 ; n3405
g3357 and n3399_not n3405 ; n3406
g3358 and n3393_not n3406 ; n3407
g3359 and n3392_not n3407 ; n3408
g3360 nor n3134 n3408 ; n3409
g3361 and n2600_not n3281 ; n3410
g3362 and n2596 n3217 ; n3411
g3363 and n2604_not n3274 ; n3412
g3364 nor n3411 n3412 ; n3413
g3365 and n3410_not n3413 ; n3414
g3366 and n2750_not n3216 ; n3415
g3367 and n3414 n3415_not ; n3416
g3368 nor n291 n3416 ; n3417
g3369 and n291 n3416 ; n3418
g3370 nor n3417 n3418 ; n3419
g3371 and n3409_not n3419 ; n3420
g3372 and n3134 n3408 ; n3421
g3373 nor n3420 n3421 ; n3422
g3374 nor n3135 n3143 ; n3423
g3375 nor n3144 n3423 ; n3424
g3376 and n3422 n3424_not ; n3425
g3377 nor n3391 n3425 ; n3426
g3378 and n3390_not n3426 ; n3427
g3379 and n3387_not n3427 ; n3428
g3380 and n3422_not n3424 ; n3429
g3381 nor n3428 n3429 ; n3430
g3382 and n2590_not n3217 ; n3431
g3383 and n2596 n3274 ; n3432
g3384 and n2593 n3281 ; n3433
g3385 nor n3432 n3433 ; n3434
g3386 and n3431_not n3434 ; n3435
g3387 and n2768 n3216 ; n3436
g3388 and n3435 n3436_not ; n3437
g3389 nor n291 n3437 ; n3438
g3390 nor n3437 n3438 ; n3439
g3391 nor n291 n3438 ; n3440
g3392 nor n3439 n3440 ; n3441
g3393 and n3430 n3441 ; n3442
g3394 nor n3156 n3442 ; n3443
g3395 and n3381_not n3443 ; n3444
g3396 nor n3430 n3441 ; n3445
g3397 nor n3444 n3445 ; n3446
g3398 nor n3160 n3171 ; n3447
g3399 and n3170 n3171_not ; n3448
g3400 nor n3447 n3448 ; n3449
g3401 and n3446 n3449 ; n3450
g3402 nor n3380 n3450 ; n3451
g3403 and n3379_not n3451 ; n3452
g3404 and n3376_not n3452 ; n3453
g3405 nor n3446 n3449 ; n3454
g3406 nor n3453 n3454 ; n3455
g3407 and n2582_not n3217 ; n3456
g3408 and n2590_not n3274 ; n3457
g3409 and n2586_not n3281 ; n3458
g3410 nor n3457 n3458 ; n3459
g3411 and n3456_not n3459 ; n3460
g3412 and n2830 n3216 ; n3461
g3413 and n3460 n3461_not ; n3462
g3414 nor n291 n3462 ; n3463
g3415 nor n3462 n3463 ; n3464
g3416 nor n291 n3463 ; n3465
g3417 nor n3464 n3465 ; n3466
g3418 and n3455 n3466 ; n3467
g3419 nor n3175 n3467 ; n3468
g3420 and n3370_not n3468 ; n3469
g3421 nor n3455 n3466 ; n3470
g3422 nor n3469 n3470 ; n3471
g3423 and n3176 n3178_not ; n3472
g3424 nor n3179 n3472 ; n3473
g3425 and n3471 n3473_not ; n3474
g3426 nor n3369 n3474 ; n3475
g3427 and n3368_not n3475 ; n3476
g3428 and n3365_not n3476 ; n3477
g3429 and n3471_not n3473 ; n3478
g3430 nor n3477 n3478 ; n3479
g3431 nor n3180 n3184 ; n3480
g3432 nor n3183 n3184 ; n3481
g3433 nor n3480 n3481 ; n3482
g3434 and n3479 n3482 ; n3483
g3435 nor n3359 n3483 ; n3484
g3436 and n3358_not n3484 ; n3485
g3437 and n3355_not n3485 ; n3486
g3438 nor n3479 n3482 ; n3487
g3439 nor n3486 n3487 ; n3488
g3440 and n3185 n3187_not ; n3489
g3441 nor n3188 n3489 ; n3490
g3442 and n3488 n3490_not ; n3491
g3443 nor n3349 n3491 ; n3492
g3444 and n3347_not n3492 ; n3493
g3445 and n3344_not n3493 ; n3494
g3446 and n3488_not n3490 ; n3495
g3447 nor n3494 n3495 ; n3496
g3448 and n3189 n3192 ; n3497
g3449 nor n3193 n3497 ; n3498
g3450 and n3496_not n3498 ; n3499
g3451 and n2566_not n3217 ; n3500
g3452 and n2575_not n3274 ; n3501
g3453 and n2562 n3281 ; n3502
g3454 nor n3501 n3502 ; n3503
g3455 and n3500_not n3503 ; n3504
g3456 and n3022 n3216 ; n3505
g3457 and n3504 n3505_not ; n3506
g3458 and n291 n3506_not ; n3507
g3459 and n291_not n3506 ; n3508
g3460 nor n3507 n3508 ; n3509
g3461 and n3499_not n3509 ; n3510
g3462 and n3496 n3498_not ; n3511
g3463 nor n3510 n3511 ; n3512
g3464 and n3194 n3197 ; n3513
g3465 nor n3198 n3513 ; n3514
g3466 nor n3512 n3514 ; n3515
g3467 and n2554_not n3217 ; n3516
g3468 and n2562 n3274 ; n3517
g3469 and n2566_not n3281 ; n3518
g3470 nor n3517 n3518 ; n3519
g3471 and n3516_not n3519 ; n3520
g3472 and n2652 n3216 ; n3521
g3473 and n3520 n3521_not ; n3522
g3474 nor n291 n3522 ; n3523
g3475 and n291 n3522 ; n3524
g3476 nor n3523 n3524 ; n3525
g3477 and n3515_not n3525 ; n3526
g3478 and n3512 n3514 ; n3527
g3479 nor n3526 n3527 ; n3528
g3480 and n3338 n3528 ; n3529
g3481 nor n3202 n3529 ; n3530
g3482 and n3325_not n3530 ; n3531
g3483 nor n3338 n3528 ; n3532
g3484 nor n3531 n3532 ; n3533
g3485 and n3310 n3324_not ; n3534
g3486 and n3323 n3324_not ; n3535
g3487 nor n3534 n3535 ; n3536
g3488 nor n3533 n3536 ; n3537
g3489 nor n3324 n3537 ; n3538
g3490 and n3208 n3308_not ; n3539
g3491 and n3307 n3308_not ; n3540
g3492 nor n3539 n3540 ; n3541
g3493 nor n3538 n3541 ; n3542
g3494 nor n3308 n3542 ; n3543
g3495 nor n3009 n3207 ; n3544
g3496 and n295 n3277 ; n3545
g3497 and n2560 n2566_not ; n3546
g3498 and n2554_not n2567 ; n3547
g3499 nor n3546 n3547 ; n3548
g3500 and n3545_not n3548 ; n3549
g3501 and n2571 n3332 ; n3550
g3502 and n3549 n3550_not ; n3551
g3503 nor n275 n3551 ; n3552
g3504 and n275 n3551 ; n3553
g3505 nor n3552 n3553 ; n3554
g3506 nor n3001 n3005 ; n3555
g3507 nor n2980 n2986 ; n3556
g3508 and n2582_not n2699 ; n3557
g3509 and n2590_not n2695 ; n3558
g3510 and n2586_not n2697 ; n3559
g3511 nor n3558 n3559 ; n3560
g3512 and n3557_not n3560 ; n3561
g3513 and n2690 n2830 ; n3562
g3514 and n3561 n3562_not ; n3563
g3515 nor n669 n3563 ; n3564
g3516 and n669 n3563 ; n3565
g3517 nor n3564 n3565 ; n3566
g3518 nor n525 n2604 ; n3567
g3519 and n2600_not n2776 ; n3568
g3520 and n2596 n2666 ; n3569
g3521 and n2593 n2668 ; n3570
g3522 nor n3569 n3570 ; n3571
g3523 and n3568_not n3571 ; n3572
g3524 and n2674 n2706_not ; n3573
g3525 and n3572 n3573_not ; n3574
g3526 nor n525 n3574 ; n3575
g3527 and n3567 n3575_not ; n3576
g3528 and n3567 n3576_not ; n3577
g3529 and n525 n3574 ; n3578
g3530 nor n3575 n3578 ; n3579
g3531 and n3576_not n3579 ; n3580
g3532 nor n3577 n3580 ; n3581
g3533 nor n2977 n3581 ; n3582
g3534 nor n2977 n3582 ; n3583
g3535 nor n3581 n3582 ; n3584
g3536 nor n3583 n3584 ; n3585
g3537 and n3566 n3585_not ; n3586
g3538 and n3566 n3586_not ; n3587
g3539 nor n3585 n3586 ; n3588
g3540 nor n3587 n3588 ; n3589
g3541 and n3556_not n3589 ; n3590
g3542 and n3556 n3589_not ; n3591
g3543 nor n3590 n3591 ; n3592
g3544 and n2562 n2802 ; n3593
g3545 and n2578 n2808 ; n3594
g3546 and n2575_not n2810 ; n3595
g3547 nor n3594 n3595 ; n3596
g3548 and n3593_not n3596 ; n3597
g3549 and n3042_not n3597 ; n3598
g3550 and n2817_not n3597 ; n3599
g3551 nor n3598 n3599 ; n3600
g3552 and n1021 n3600_not ; n3601
g3553 and n1021_not n3600 ; n3602
g3554 nor n3601 n3602 ; n3603
g3555 and n3592_not n3603 ; n3604
g3556 and n3592 n3603_not ; n3605
g3557 nor n3604 n3605 ; n3606
g3558 and n3555_not n3606 ; n3607
g3559 and n3555 n3606_not ; n3608
g3560 nor n3607 n3608 ; n3609
g3561 and n3554 n3609 ; n3610
g3562 nor n3554 n3609 ; n3611
g3563 nor n3610 n3611 ; n3612
g3564 and n3544_not n3612 ; n3613
g3565 and n3544 n3612_not ; n3614
g3566 nor n3613 n3614 ; n3615
g3567 and n348_not n502 ; n3616
g3568 and n148_not n3616 ; n3617
g3569 and n514 n3617 ; n3618
g3570 and n485 n3618 ; n3619
g3571 and n414 n3619 ; n3620
g3572 and n404 n3620 ; n3621
g3573 and n188_not n3621 ; n3622
g3574 and n219_not n3622 ; n3623
g3575 and n224_not n3623 ; n3624
g3576 and n3258 n3269 ; n3625
g3577 nor n3624 n3625 ; n3626
g3578 and n3624 n3625 ; n3627
g3579 nor n3626 n3627 ; n3628
g3580 and n3217 n3628_not ; n3629
g3581 and n3274 n3280_not ; n3630
g3582 and n3272 n3281 ; n3631
g3583 nor n3630 n3631 ; n3632
g3584 and n3629_not n3632 ; n3633
g3585 and n3216_not n3633 ; n3634
g3586 nor n3298 n3300 ; n3635
g3587 and n3272_not n3628 ; n3636
g3588 and n3272 n3628_not ; n3637
g3589 nor n3636 n3637 ; n3638
g3590 and n3635_not n3638 ; n3639
g3591 and n3635 n3638_not ; n3640
g3592 nor n3639 n3640 ; n3641
g3593 and n3633 n3641_not ; n3642
g3594 nor n3634 n3642 ; n3643
g3595 and n291 n3643_not ; n3644
g3596 and n291_not n3643 ; n3645
g3597 nor n3644 n3645 ; n3646
g3598 and n3615 n3646 ; n3647
g3599 nor n3615 n3646 ; n3648
g3600 nor n3647 n3648 ; n3649
g3601 and n3543_not n3649 ; n3650
g3602 and n3543 n3649_not ; n3651
g3603 nor n3650 n3651 ; n3652
g3604 and n271_not n3652 ; n3653
g3605 nor n114 n506 ; n3654
g3606 and n736_not n3654 ; n3655
g3607 and n296_not n3655 ; n3656
g3608 and n154_not n3656 ; n3657
g3609 and n806 n3657 ; n3658
g3610 and n139_not n3658 ; n3659
g3611 and n150_not n3659 ; n3660
g3612 and n186_not n3660 ; n3661
g3613 and n313_not n3661 ; n3662
g3614 and n133_not n3662 ; n3663
g3615 and n359_not n3663 ; n3664
g3616 and n142_not n3664 ; n3665
g3617 and n106_not n3665 ; n3666
g3618 and n372 n505 ; n3667
g3619 and n1134 n3667 ; n3668
g3620 and n217_not n3668 ; n3669
g3621 and n255_not n3669 ; n3670
g3622 and n495_not n3670 ; n3671
g3623 and n553_not n3671 ; n3672
g3624 and n445_not n3672 ; n3673
g3625 and n471_not n3673 ; n3674
g3626 and n215_not n3674 ; n3675
g3627 and n789 n3675 ; n3676
g3628 and n417_not n3676 ; n3677
g3629 and n298_not n3677 ; n3678
g3630 and n2454 n3678 ; n3679
g3631 and n3666 n3679 ; n3680
g3632 and n980 n3680 ; n3681
g3633 and n137_not n3681 ; n3682
g3634 and n254_not n3682 ; n3683
g3635 and n327_not n3683 ; n3684
g3636 and n446_not n3684 ; n3685
g3637 and n146_not n3685 ; n3686
g3638 and n297_not n3686 ; n3687
g3639 and n335_not n3687 ; n3688
g3640 and n470_not n3688 ; n3689
g3641 and n342_not n3689 ; n3690
g3642 and n3538 n3540_not ; n3691
g3643 and n3539_not n3691 ; n3692
g3644 nor n3542 n3692 ; n3693
g3645 and n397 n2278 ; n3694
g3646 and n2303 n3694 ; n3695
g3647 and n144_not n3695 ; n3696
g3648 and n503_not n3696 ; n3697
g3649 and n356_not n3697 ; n3698
g3650 and n477_not n3698 ; n3699
g3651 and n341 n813 ; n3700
g3652 and n137_not n3700 ; n3701
g3653 and n155_not n3701 ; n3702
g3654 and n460 n2422 ; n3703
g3655 and n2433 n3703 ; n3704
g3656 and n344 n3704 ; n3705
g3657 and n3702 n3705 ; n3706
g3658 and n3699 n3706 ; n3707
g3659 and n2364 n3707 ; n3708
g3660 and n415_not n3708 ; n3709
g3661 and n150_not n3709 ; n3710
g3662 and n317_not n3710 ; n3711
g3663 and n219_not n3711 ; n3712
g3664 and n174_not n3712 ; n3713
g3665 and n218_not n3713 ; n3714
g3666 and n302_not n3714 ; n3715
g3667 and n3533 n3536 ; n3716
g3668 nor n3537 n3716 ; n3717
g3669 and n3715_not n3717 ; n3718
g3670 nor n3693 n3718 ; n3719
g3671 nor n3690 n3719 ; n3720
g3672 and n3693 n3718 ; n3721
g3673 nor n3720 n3721 ; n3722
g3674 nor n271 n3653 ; n3723
g3675 and n3652 n3653_not ; n3724
g3676 nor n3723 n3724 ; n3725
g3677 nor n3722 n3725 ; n3726
g3678 nor n3653 n3726 ; n3727
g3679 and n239 n590 ; n3728
g3680 and n350_not n3728 ; n3729
g3681 and n123_not n3729 ; n3730
g3682 and n313_not n3730 ; n3731
g3683 and n207_not n3731 ; n3732
g3684 and n445_not n3732 ; n3733
g3685 and n469_not n3733 ; n3734
g3686 and n353 n468_not ; n3735
g3687 and n334 n3735 ; n3736
g3688 and n1162 n3736 ; n3737
g3689 and n3734 n3737 ; n3738
g3690 and n2418 n3738 ; n3739
g3691 and n222_not n3739 ; n3740
g3692 and n317_not n3740 ; n3741
g3693 and n177_not n3741 ; n3742
g3694 and n218_not n3742 ; n3743
g3695 and n554_not n3743 ; n3744
g3696 and n211_not n3744 ; n3745
g3697 and n132_not n3745 ; n3746
g3698 and n223_not n3746 ; n3747
g3699 and n3627_not n3747 ; n3748
g3700 and n3627 n3747_not ; n3749
g3701 nor n3748 n3749 ; n3750
g3702 and n3217 n3750 ; n3751
g3703 and n3272 n3274 ; n3752
g3704 and n3281 n3628_not ; n3753
g3705 nor n3752 n3753 ; n3754
g3706 and n3751_not n3754 ; n3755
g3707 nor n3637 n3639 ; n3756
g3708 and n3628 n3750_not ; n3757
g3709 and n3628_not n3750 ; n3758
g3710 nor n3757 n3758 ; n3759
g3711 and n3756_not n3759 ; n3760
g3712 and n3756 n3759_not ; n3761
g3713 nor n3760 n3761 ; n3762
g3714 and n3216 n3762 ; n3763
g3715 and n3755 n3763_not ; n3764
g3716 nor n291 n3764 ; n3765
g3717 nor n3764 n3765 ; n3766
g3718 nor n291 n3765 ; n3767
g3719 nor n3766 n3767 ; n3768
g3720 nor n3610 n3613 ; n3769
g3721 and n2566_not n2802 ; n3770
g3722 and n2575_not n2808 ; n3771
g3723 and n2562 n2810 ; n3772
g3724 nor n3771 n3772 ; n3773
g3725 and n3770_not n3773 ; n3774
g3726 and n2817 n3022 ; n3775
g3727 and n3774 n3775_not ; n3776
g3728 nor n1021 n3776 ; n3777
g3729 nor n3776 n3777 ; n3778
g3730 nor n1021 n3777 ; n3779
g3731 nor n3778 n3779 ; n3780
g3732 nor n3556 n3589 ; n3781
g3733 nor n3586 n3781 ; n3782
g3734 nor n3576 n3582 ; n3783
g3735 and n2590_not n2668 ; n3784
g3736 and n2596 n2776 ; n3785
g3737 and n2593 n2666 ; n3786
g3738 nor n3785 n3786 ; n3787
g3739 and n3784_not n3787 ; n3788
g3740 and n2674 n2768 ; n3789
g3741 and n3788 n3789_not ; n3790
g3742 and n525_not n2600 ; n3791
g3743 and n3790_not n3791 ; n3792
g3744 and n3790 n3791_not ; n3793
g3745 nor n3792 n3793 ; n3794
g3746 and n3783_not n3794 ; n3795
g3747 and n3783 n3794_not ; n3796
g3748 nor n3795 n3796 ; n3797
g3749 and n2578 n2699 ; n3798
g3750 and n2586_not n2695 ; n3799
g3751 and n2582_not n2697 ; n3800
g3752 nor n3799 n3800 ; n3801
g3753 and n3798_not n3801 ; n3802
g3754 and n2690_not n3802 ; n3803
g3755 and n2815_not n3802 ; n3804
g3756 nor n3803 n3804 ; n3805
g3757 and n669 n3805_not ; n3806
g3758 and n669_not n3805 ; n3807
g3759 nor n3806 n3807 ; n3808
g3760 and n3797 n3808 ; n3809
g3761 and n3797 n3809_not ; n3810
g3762 and n3808 n3809_not ; n3811
g3763 nor n3810 n3811 ; n3812
g3764 nor n3782 n3812 ; n3813
g3765 nor n3782 n3813 ; n3814
g3766 nor n3812 n3813 ; n3815
g3767 nor n3814 n3815 ; n3816
g3768 nor n3780 n3816 ; n3817
g3769 nor n3780 n3817 ; n3818
g3770 nor n3816 n3817 ; n3819
g3771 nor n3818 n3819 ; n3820
g3772 nor n3604 n3607 ; n3821
g3773 and n3820 n3821 ; n3822
g3774 nor n3820 n3821 ; n3823
g3775 nor n3822 n3823 ; n3824
g3776 and n295 n3280_not ; n3825
g3777 and n2554_not n2560 ; n3826
g3778 and n2567 n3277 ; n3827
g3779 nor n3826 n3827 ; n3828
g3780 and n3825_not n3828 ; n3829
g3781 and n2571_not n3829 ; n3830
g3782 and n3318_not n3829 ; n3831
g3783 nor n3830 n3831 ; n3832
g3784 and n275 n3832_not ; n3833
g3785 and n275_not n3832 ; n3834
g3786 nor n3833 n3834 ; n3835
g3787 and n3824 n3835 ; n3836
g3788 and n3824 n3836_not ; n3837
g3789 and n3835 n3836_not ; n3838
g3790 nor n3837 n3838 ; n3839
g3791 nor n3769 n3839 ; n3840
g3792 nor n3769 n3840 ; n3841
g3793 nor n3839 n3840 ; n3842
g3794 nor n3841 n3842 ; n3843
g3795 nor n3768 n3843 ; n3844
g3796 nor n3768 n3844 ; n3845
g3797 nor n3843 n3844 ; n3846
g3798 nor n3845 n3846 ; n3847
g3799 nor n3647 n3650 ; n3848
g3800 and n3847 n3848 ; n3849
g3801 nor n3847 n3848 ; n3850
g3802 nor n3849 n3850 ; n3851
g3803 and n239 n1093 ; n3852
g3804 and n806 n3852 ; n3853
g3805 and n1459 n3853 ; n3854
g3806 and n2311 n3854 ; n3855
g3807 and n643 n3855 ; n3856
g3808 and n623 n3856 ; n3857
g3809 and n210 n3857 ; n3858
g3810 and n255_not n3858 ; n3859
g3811 and n148_not n3859 ; n3860
g3812 and n345_not n3860 ; n3861
g3813 and n3851_not n3861 ; n3862
g3814 and n3851 n3861_not ; n3863
g3815 nor n3862 n3863 ; n3864
g3816 and n3727_not n3864 ; n3865
g3817 and n3727 n3864_not ; n3866
g3818 nor n3865 n3866 ; n3867
g3819 nor n3722 n3726 ; n3868
g3820 nor n3725 n3726 ; n3869
g3821 nor n3868 n3869 ; n3870
g3822 and n3867 n3870_not ; n3871
g3823 and n3867 n3871_not ; n3872
g3824 nor n3870 n3871 ; n3873
g3825 or n3872 n3873 ; sin[0]
g3826 nor n3863 n3865 ; n3875
g3827 and n3627 n3747 ; n3876
g3828 and n236 n2433 ; n3877
g3829 and n457 n3877 ; n3878
g3830 and n753 n3878 ; n3879
g3831 and n169_not n3879 ; n3880
g3832 and n118_not n3880 ; n3881
g3833 and n166_not n3881 ; n3882
g3834 and n168_not n3882 ; n3883
g3835 and n316 n555 ; n3884
g3836 and n815 n3884 ; n3885
g3837 and n1476 n3885 ; n3886
g3838 and n3883 n3886 ; n3887
g3839 and n2432 n3887 ; n3888
g3840 and n976 n3888 ; n3889
g3841 and n495_not n3889 ; n3890
g3842 and n470_not n3890 ; n3891
g3843 and n367_not n3891 ; n3892
g3844 and n326_not n3892 ; n3893
g3845 and n3876_not n3893 ; n3894
g3846 and n3876 n3893_not ; n3895
g3847 nor n3894 n3895 ; n3896
g3848 and n3217 n3896 ; n3897
g3849 and n3274 n3628_not ; n3898
g3850 and n3281 n3750 ; n3899
g3851 nor n3898 n3899 ; n3900
g3852 and n3897_not n3900 ; n3901
g3853 nor n3758 n3760 ; n3902
g3854 nor n3750 n3896 ; n3903
g3855 and n3750 n3896 ; n3904
g3856 nor n3903 n3904 ; n3905
g3857 and n3902_not n3905 ; n3906
g3858 and n3902 n3905_not ; n3907
g3859 nor n3906 n3907 ; n3908
g3860 and n3216 n3908 ; n3909
g3861 and n3901 n3909_not ; n3910
g3862 nor n291 n3910 ; n3911
g3863 nor n3910 n3911 ; n3912
g3864 nor n291 n3911 ; n3913
g3865 nor n3912 n3913 ; n3914
g3866 nor n3836 n3840 ; n3915
g3867 and n2554_not n2802 ; n3916
g3868 and n2562 n2808 ; n3917
g3869 and n2566_not n2810 ; n3918
g3870 nor n3917 n3918 ; n3919
g3871 and n3916_not n3919 ; n3920
g3872 and n2652 n2817 ; n3921
g3873 and n3920 n3921_not ; n3922
g3874 nor n1021 n3922 ; n3923
g3875 nor n3922 n3923 ; n3924
g3876 nor n1021 n3923 ; n3925
g3877 nor n3924 n3925 ; n3926
g3878 nor n3809 n3813 ; n3927
g3879 nor n525 n2600 ; n3928
g3880 and n3790 n3928 ; n3929
g3881 nor n3795 n3929 ; n3930
g3882 and n2586_not n2668 ; n3931
g3883 and n2593 n2776 ; n3932
g3884 and n2590_not n2666 ; n3933
g3885 nor n3932 n3933 ; n3934
g3886 and n3931_not n3934 ; n3935
g3887 and n2674 n2849 ; n3936
g3888 and n3935 n3936_not ; n3937
g3889 nor n525 n2596 ; n3938
g3890 and n3937_not n3938 ; n3939
g3891 and n3937 n3938_not ; n3940
g3892 nor n3939 n3940 ; n3941
g3893 and n3930_not n3941 ; n3942
g3894 nor n3930 n3942 ; n3943
g3895 and n3941 n3942_not ; n3944
g3896 nor n3943 n3944 ; n3945
g3897 and n2575_not n2699 ; n3946
g3898 and n2582_not n2695 ; n3947
g3899 and n2578 n2697 ; n3948
g3900 nor n3947 n3948 ; n3949
g3901 and n3946_not n3949 ; n3950
g3902 and n2690_not n3950 ; n3951
g3903 and n2989_not n3950 ; n3952
g3904 nor n3951 n3952 ; n3953
g3905 and n669 n3953_not ; n3954
g3906 and n669_not n3953 ; n3955
g3907 nor n3954 n3955 ; n3956
g3908 and n3945_not n3956 ; n3957
g3909 nor n3945 n3957 ; n3958
g3910 and n3956 n3957_not ; n3959
g3911 nor n3958 n3959 ; n3960
g3912 nor n3927 n3960 ; n3961
g3913 nor n3927 n3961 ; n3962
g3914 nor n3960 n3961 ; n3963
g3915 nor n3962 n3963 ; n3964
g3916 nor n3926 n3964 ; n3965
g3917 nor n3926 n3965 ; n3966
g3918 nor n3964 n3965 ; n3967
g3919 nor n3966 n3967 ; n3968
g3920 nor n3817 n3823 ; n3969
g3921 and n3968 n3969 ; n3970
g3922 nor n3968 n3969 ; n3971
g3923 nor n3970 n3971 ; n3972
g3924 and n295 n3272 ; n3973
g3925 and n2560 n3277 ; n3974
g3926 and n2567 n3280_not ; n3975
g3927 nor n3974 n3975 ; n3976
g3928 and n3973_not n3976 ; n3977
g3929 and n2571_not n3977 ; n3978
g3930 and n3302_not n3977 ; n3979
g3931 nor n3978 n3979 ; n3980
g3932 and n275 n3980_not ; n3981
g3933 and n275_not n3980 ; n3982
g3934 nor n3981 n3982 ; n3983
g3935 and n3972 n3983 ; n3984
g3936 and n3972 n3984_not ; n3985
g3937 and n3983 n3984_not ; n3986
g3938 nor n3985 n3986 ; n3987
g3939 nor n3915 n3987 ; n3988
g3940 nor n3915 n3988 ; n3989
g3941 nor n3987 n3988 ; n3990
g3942 nor n3989 n3990 ; n3991
g3943 nor n3914 n3991 ; n3992
g3944 nor n3914 n3992 ; n3993
g3945 nor n3991 n3992 ; n3994
g3946 nor n3993 n3994 ; n3995
g3947 nor n3844 n3850 ; n3996
g3948 and n3995 n3996 ; n3997
g3949 nor n3995 n3996 ; n3998
g3950 nor n3997 n3998 ; n3999
g3951 nor n140 n405 ; n4000
g3952 and n361_not n4000 ; n4001
g3953 and n258_not n4001 ; n4002
g3954 and n637 n2340 ; n4003
g3955 and n2276 n4003 ; n4004
g3956 and n249 n4004 ; n4005
g3957 and n753 n4005 ; n4006
g3958 and n4002 n4006 ; n4007
g3959 and n210 n4007 ; n4008
g3960 and n3231 n4008 ; n4009
g3961 and n175_not n4009 ; n4010
g3962 and n155_not n4010 ; n4011
g3963 and n327_not n4011 ; n4012
g3964 and n191_not n4012 ; n4013
g3965 and n118_not n4013 ; n4014
g3966 and n445_not n4014 ; n4015
g3967 and n3999_not n4015 ; n4016
g3968 and n3999 n4015_not ; n4017
g3969 nor n4016 n4017 ; n4018
g3970 and n3875_not n4018 ; n4019
g3971 and n3875 n4018_not ; n4020
g3972 nor n4019 n4020 ; n4021
g3973 and n3871 n4021 ; n4022
g3974 nor n3871 n4021 ; n4023
g3975 nor n4022 n4023 ; n4024
g3976 and a[22] a[23]_not ; n4025
g3977 and a[22]_not a[23] ; n4026
g3978 nor n4025 n4026 ; n4027
g3979 and sin[0] n4027_not ; n4028
g3980 and n4024_not n4028 ; n4029
g3981 and n4024 n4028_not ; n4030
g3982 or n4029 n4030 ; sin[1]
g3983 nor n4017 n4019 ; n4032
g3984 and n346 n408_not ; n4033
g3985 and n129_not n4033 ; n4034
g3986 and n228_not n4034 ; n4035
g3987 and n142_not n4035 ; n4036
g3988 and n132_not n4036 ; n4037
g3989 and n416 n608 ; n4038
g3990 and n805 n4038 ; n4039
g3991 and n4037 n4039 ; n4040
g3992 and n3699 n4040 ; n4041
g3993 and n313_not n4041 ; n4042
g3994 and n458_not n4042 ; n4043
g3995 and n504_not n4043 ; n4044
g3996 and n298_not n4044 ; n4045
g3997 and n146_not n4045 ; n4046
g3998 and n506_not n4046 ; n4047
g3999 and n326_not n4047 ; n4048
g4000 nor n3992 n3998 ; n4049
g4001 and n3274 n3750 ; n4050
g4002 and n3281 n3896 ; n4051
g4003 nor n4050 n4051 ; n4052
g4004 nor n3750 n3906 ; n4053
g4005 and n3896 n4053_not ; n4054
g4006 nor n3896 n3906 ; n4055
g4007 nor n4054 n4055 ; n4056
g4008 and n3216 n4056 ; n4057
g4009 and n4052 n4057_not ; n4058
g4010 nor n291 n4058 ; n4059
g4011 nor n4058 n4059 ; n4060
g4012 nor n291 n4059 ; n4061
g4013 nor n4060 n4061 ; n4062
g4014 nor n3984 n3988 ; n4063
g4015 and n2802 n3277 ; n4064
g4016 and n2566_not n2808 ; n4065
g4017 and n2554_not n2810 ; n4066
g4018 nor n4065 n4066 ; n4067
g4019 and n4064_not n4067 ; n4068
g4020 and n2817 n3332 ; n4069
g4021 and n4068 n4069_not ; n4070
g4022 nor n1021 n4070 ; n4071
g4023 nor n4070 n4071 ; n4072
g4024 nor n1021 n4071 ; n4073
g4025 nor n4072 n4073 ; n4074
g4026 nor n3957 n3961 ; n4075
g4027 and n525_not n3937 ; n4076
g4028 and n2596 n4076 ; n4077
g4029 nor n3942 n4077 ; n4078
g4030 and n2582_not n2668 ; n4079
g4031 and n2590_not n2776 ; n4080
g4032 and n2586_not n2666 ; n4081
g4033 nor n4080 n4081 ; n4082
g4034 and n4079_not n4082 ; n4083
g4035 and n2674 n2830 ; n4084
g4036 and n4083 n4084_not ; n4085
g4037 nor n525 n2593 ; n4086
g4038 and n4085_not n4086 ; n4087
g4039 and n4085 n4086_not ; n4088
g4040 nor n4087 n4088 ; n4089
g4041 and n4078_not n4089 ; n4090
g4042 nor n4078 n4090 ; n4091
g4043 and n4089 n4090_not ; n4092
g4044 nor n4091 n4092 ; n4093
g4045 and n2562 n2699 ; n4094
g4046 and n2578 n2695 ; n4095
g4047 and n2575_not n2697 ; n4096
g4048 nor n4095 n4096 ; n4097
g4049 and n4094_not n4097 ; n4098
g4050 and n2690_not n4098 ; n4099
g4051 and n3042_not n4098 ; n4100
g4052 nor n4099 n4100 ; n4101
g4053 and n669 n4101_not ; n4102
g4054 and n669_not n4101 ; n4103
g4055 nor n4102 n4103 ; n4104
g4056 and n4093_not n4104 ; n4105
g4057 nor n4093 n4105 ; n4106
g4058 and n4104 n4105_not ; n4107
g4059 nor n4106 n4107 ; n4108
g4060 nor n4075 n4108 ; n4109
g4061 nor n4075 n4109 ; n4110
g4062 nor n4108 n4109 ; n4111
g4063 nor n4110 n4111 ; n4112
g4064 nor n4074 n4112 ; n4113
g4065 nor n4074 n4113 ; n4114
g4066 nor n4112 n4113 ; n4115
g4067 nor n4114 n4115 ; n4116
g4068 nor n3965 n3971 ; n4117
g4069 and n4116 n4117 ; n4118
g4070 nor n4116 n4117 ; n4119
g4071 nor n4118 n4119 ; n4120
g4072 and n295 n3628_not ; n4121
g4073 and n2560 n3280_not ; n4122
g4074 and n2567 n3272 ; n4123
g4075 nor n4122 n4123 ; n4124
g4076 and n4121_not n4124 ; n4125
g4077 and n2571_not n4125 ; n4126
g4078 and n3641_not n4125 ; n4127
g4079 nor n4126 n4127 ; n4128
g4080 and n275 n4128_not ; n4129
g4081 and n275_not n4128 ; n4130
g4082 nor n4129 n4130 ; n4131
g4083 and n4120 n4131 ; n4132
g4084 and n4120 n4132_not ; n4133
g4085 and n4131 n4132_not ; n4134
g4086 nor n4133 n4134 ; n4135
g4087 nor n4063 n4135 ; n4136
g4088 nor n4063 n4136 ; n4137
g4089 nor n4135 n4136 ; n4138
g4090 nor n4137 n4138 ; n4139
g4091 nor n4062 n4139 ; n4140
g4092 nor n4062 n4140 ; n4141
g4093 nor n4139 n4140 ; n4142
g4094 nor n4141 n4142 ; n4143
g4095 and n4049_not n4143 ; n4144
g4096 and n4049 n4143_not ; n4145
g4097 nor n4144 n4145 ; n4146
g4098 nor n4048 n4146 ; n4147
g4099 and n4048 n4146 ; n4148
g4100 nor n4032 n4148 ; n4149
g4101 and n4147_not n4149 ; n4150
g4102 nor n4032 n4150 ; n4151
g4103 nor n4147 n4150 ; n4152
g4104 and n4148_not n4152 ; n4153
g4105 nor n4151 n4153 ; n4154
g4106 and n4022_not n4154 ; n4155
g4107 and n4022 n4154_not ; n4156
g4108 nor n4155 n4156 ; n4157
g4109 nor sin[0] n4024 ; n4158
g4110 nor n4027 n4158 ; n4159
g4111 and n4157_not n4159 ; n4160
g4112 and n4157 n4159_not ; n4161
g4113 or n4160 n4161 ; sin[2]
g4114 and n2340 n3657 ; n4163
g4115 and n397 n4163 ; n4164
g4116 and n946 n4164 ; n4165
g4117 and n2196 n4165 ; n4166
g4118 and n1468 n4166 ; n4167
g4119 and n735 n4167 ; n4168
g4120 and n355 n4168 ; n4169
g4121 and n317_not n4169 ; n4170
g4122 and n175_not n4170 ; n4171
g4123 and n370_not n4171 ; n4172
g4124 and n111_not n4172 ; n4173
g4125 and n258_not n4173 ; n4174
g4126 and n238_not n4174 ; n4175
g4127 nor n4049 n4143 ; n4176
g4128 nor n4140 n4176 ; n4177
g4129 nor n4132 n4136 ; n4178
g4130 and n3274 n3896 ; n4179
g4131 and n3216 n4054 ; n4180
g4132 nor n4179 n4180 ; n4181
g4133 nor n291 n4181 ; n4182
g4134 nor n4181 n4182 ; n4183
g4135 nor n291 n4182 ; n4184
g4136 nor n4183 n4184 ; n4185
g4137 and n2802 n3280_not ; n4186
g4138 and n2554_not n2808 ; n4187
g4139 and n2810 n3277 ; n4188
g4140 nor n4187 n4188 ; n4189
g4141 and n4186_not n4189 ; n4190
g4142 and n2817 n3318 ; n4191
g4143 and n4190 n4191_not ; n4192
g4144 nor n1021 n4192 ; n4193
g4145 nor n4192 n4193 ; n4194
g4146 nor n1021 n4193 ; n4195
g4147 nor n4194 n4195 ; n4196
g4148 nor n4105 n4109 ; n4197
g4149 and n525_not n4085 ; n4198
g4150 and n2593 n4198 ; n4199
g4151 nor n4090 n4199 ; n4200
g4152 and n2578 n2668 ; n4201
g4153 and n2586_not n2776 ; n4202
g4154 and n2582_not n2666 ; n4203
g4155 nor n4202 n4203 ; n4204
g4156 and n4201_not n4204 ; n4205
g4157 and n2674 n2815 ; n4206
g4158 and n4205 n4206_not ; n4207
g4159 and n525_not n2590 ; n4208
g4160 and n4207_not n4208 ; n4209
g4161 and n4207 n4208_not ; n4210
g4162 nor n4209 n4210 ; n4211
g4163 and n4200_not n4211 ; n4212
g4164 nor n4200 n4212 ; n4213
g4165 and n4211 n4212_not ; n4214
g4166 nor n4213 n4214 ; n4215
g4167 and n2566_not n2699 ; n4216
g4168 and n2575_not n2695 ; n4217
g4169 and n2562 n2697 ; n4218
g4170 nor n4217 n4218 ; n4219
g4171 and n4216_not n4219 ; n4220
g4172 and n2690_not n4220 ; n4221
g4173 and n3022_not n4220 ; n4222
g4174 nor n4221 n4222 ; n4223
g4175 and n669 n4223_not ; n4224
g4176 and n669_not n4223 ; n4225
g4177 nor n4224 n4225 ; n4226
g4178 and n4215_not n4226 ; n4227
g4179 and n4215 n4226_not ; n4228
g4180 nor n4227 n4228 ; n4229
g4181 and n4197_not n4229 ; n4230
g4182 and n4197 n4229_not ; n4231
g4183 nor n4230 n4231 ; n4232
g4184 and n4196_not n4232 ; n4233
g4185 nor n4196 n4233 ; n4234
g4186 and n4232 n4233_not ; n4235
g4187 nor n4234 n4235 ; n4236
g4188 nor n4113 n4119 ; n4237
g4189 and n4236 n4237 ; n4238
g4190 nor n4236 n4237 ; n4239
g4191 nor n4238 n4239 ; n4240
g4192 and n295 n3750 ; n4241
g4193 and n2560 n3272 ; n4242
g4194 and n2567 n3628_not ; n4243
g4195 nor n4242 n4243 ; n4244
g4196 and n4241_not n4244 ; n4245
g4197 and n2571_not n4245 ; n4246
g4198 and n3762_not n4245 ; n4247
g4199 nor n4246 n4247 ; n4248
g4200 and n275 n4248_not ; n4249
g4201 and n275_not n4248 ; n4250
g4202 nor n4249 n4250 ; n4251
g4203 and n4240 n4251 ; n4252
g4204 nor n4240 n4251 ; n4253
g4205 nor n4252 n4253 ; n4254
g4206 and n4185_not n4254 ; n4255
g4207 and n4185 n4254_not ; n4256
g4208 nor n4255 n4256 ; n4257
g4209 and n4178_not n4257 ; n4258
g4210 and n4178 n4257_not ; n4259
g4211 nor n4258 n4259 ; n4260
g4212 and n4177_not n4260 ; n4261
g4213 and n4177 n4260_not ; n4262
g4214 nor n4261 n4262 ; n4263
g4215 and n4175_not n4263 ; n4264
g4216 nor n4175 n4264 ; n4265
g4217 and n4263 n4264_not ; n4266
g4218 nor n4265 n4266 ; n4267
g4219 nor n4152 n4267 ; n4268
g4220 and n4152 n4266_not ; n4269
g4221 and n4265_not n4269 ; n4270
g4222 nor n4268 n4270 ; n4271
g4223 and n4156 n4271 ; n4272
g4224 and n4271 n4272_not ; n4273
g4225 and n4156 n4272_not ; n4274
g4226 nor n4273 n4274 ; n4275
g4227 and n4157_not n4158 ; n4276
g4228 nor n4027 n4276 ; n4277
g4229 and n4275_not n4277 ; n4278
g4230 and n4275 n4277_not ; n4279
g4231 nor n4278 n4279 ; sin[3]
g4232 nor n4264 n4268 ; n4281
g4233 and n346 n496 ; n4282
g4234 and n301 n4282 ; n4283
g4235 and n2464 n4283 ; n4284
g4236 and n975 n4284 ; n4285
g4237 and n752 n4285 ; n4286
g4238 and n644 n4286 ; n4287
g4239 and n2418 n4287 ; n4288
g4240 and n178_not n4288 ; n4289
g4241 and n194_not n4289 ; n4290
g4242 and n589_not n4290 ; n4291
g4243 nor n4258 n4261 ; n4292
g4244 nor n4252 n4255 ; n4293
g4245 nor n4233 n4239 ; n4294
g4246 nor n4227 n4230 ; n4295
g4247 and n2575_not n2668 ; n4296
g4248 and n2582_not n2776 ; n4297
g4249 and n2578 n2666 ; n4298
g4250 nor n4297 n4298 ; n4299
g4251 and n4296_not n4299 ; n4300
g4252 and n2674 n2989 ; n4301
g4253 and n4300 n4301_not ; n4302
g4254 nor n525 n4302 ; n4303
g4255 nor n4302 n4303 ; n4304
g4256 nor n525 n4303 ; n4305
g4257 nor n4304 n4305 ; n4306
g4258 nor n291 n525 ; n4307
g4259 and n2586_not n4307 ; n4308
g4260 nor n291 n4308 ; n4309
g4261 nor n2586 n4308 ; n4310
g4262 and n525_not n4310 ; n4311
g4263 nor n4309 n4311 ; n4312
g4264 nor n4306 n4312 ; n4313
g4265 nor n4306 n4313 ; n4314
g4266 nor n4312 n4313 ; n4315
g4267 nor n4314 n4315 ; n4316
g4268 nor n525 n2590 ; n4317
g4269 and n4207 n4317 ; n4318
g4270 nor n4212 n4318 ; n4319
g4271 and n4316 n4319_not ; n4320
g4272 and n4316_not n4319 ; n4321
g4273 nor n4320 n4321 ; n4322
g4274 and n2554_not n2699 ; n4323
g4275 and n2562 n2695 ; n4324
g4276 and n2566_not n2697 ; n4325
g4277 nor n4324 n4325 ; n4326
g4278 and n4323_not n4326 ; n4327
g4279 and n2652 n2690 ; n4328
g4280 and n4327 n4328_not ; n4329
g4281 nor n669 n4329 ; n4330
g4282 and n669 n4329 ; n4331
g4283 nor n4330 n4331 ; n4332
g4284 and n4322_not n4332 ; n4333
g4285 nor n4322 n4333 ; n4334
g4286 and n4332 n4333_not ; n4335
g4287 nor n4334 n4335 ; n4336
g4288 and n4295_not n4336 ; n4337
g4289 and n4295 n4336_not ; n4338
g4290 nor n4337 n4338 ; n4339
g4291 and n2802 n3272 ; n4340
g4292 and n2808 n3277 ; n4341
g4293 and n2810 n3280_not ; n4342
g4294 nor n4341 n4342 ; n4343
g4295 and n4340_not n4343 ; n4344
g4296 and n2817 n3302 ; n4345
g4297 and n4344 n4345_not ; n4346
g4298 nor n1021 n4346 ; n4347
g4299 nor n1021 n4347 ; n4348
g4300 nor n4346 n4347 ; n4349
g4301 nor n4348 n4349 ; n4350
g4302 nor n4339 n4350 ; n4351
g4303 and n4339 n4350 ; n4352
g4304 nor n4351 n4352 ; n4353
g4305 and n4294_not n4353 ; n4354
g4306 and n4294 n4353_not ; n4355
g4307 nor n4354 n4355 ; n4356
g4308 and n295 n3896 ; n4357
g4309 and n2560 n3628_not ; n4358
g4310 and n2567 n3750 ; n4359
g4311 nor n4358 n4359 ; n4360
g4312 and n4357_not n4360 ; n4361
g4313 and n2571 n3908 ; n4362
g4314 and n4361 n4362_not ; n4363
g4315 nor n275 n4363 ; n4364
g4316 and n275 n4363 ; n4365
g4317 nor n4364 n4365 ; n4366
g4318 and n4356 n4366 ; n4367
g4319 nor n4356 n4366 ; n4368
g4320 nor n4367 n4368 ; n4369
g4321 and n4293_not n4369 ; n4370
g4322 and n4293 n4369_not ; n4371
g4323 nor n4370 n4371 ; n4372
g4324 and n4292 n4372_not ; n4373
g4325 and n4292_not n4372 ; n4374
g4326 nor n4373 n4374 ; n4375
g4327 and n4291 n4375_not ; n4376
g4328 and n4291_not n4375 ; n4377
g4329 nor n4376 n4377 ; n4378
g4330 and n4281_not n4378 ; n4379
g4331 and n4281 n4378_not ; n4380
g4332 nor n4379 n4380 ; n4381
g4333 nor n4272 n4381 ; n4382
g4334 and n4272 n4381 ; n4383
g4335 nor n4382 n4383 ; n4384
g4336 and n4275 n4276 ; n4385
g4337 nor n4027 n4385 ; n4386
g4338 and n4384_not n4386 ; n4387
g4339 and n4384 n4386_not ; n4388
g4340 or n4387 n4388 ; sin[4]
g4341 nor n4377 n4379 ; n4390
g4342 nor n317 n359 ; n4391
g4343 and n472_not n4391 ; n4392
g4344 and n189 n807 ; n4393
g4345 and n4392 n4393 ; n4394
g4346 and n2317 n4394 ; n4395
g4347 and n314 n4395 ; n4396
g4348 and n3883 n4396 ; n4397
g4349 and n3243 n4397 ; n4398
g4350 and n4002 n4398 ; n4399
g4351 and n369 n4399 ; n4400
g4352 and n178_not n4400 ; n4401
g4353 and n417_not n4401 ; n4402
g4354 and n299_not n4402 ; n4403
g4355 and n237_not n4403 ; n4404
g4356 nor n4370 n4374 ; n4405
g4357 nor n4354 n4367 ; n4406
g4358 nor n4295 n4336 ; n4407
g4359 nor n4351 n4407 ; n4408
g4360 and n2802 n3628_not ; n4409
g4361 and n2808 n3280_not ; n4410
g4362 and n2810 n3272 ; n4411
g4363 nor n4410 n4411 ; n4412
g4364 and n4409_not n4412 ; n4413
g4365 and n2817 n3641 ; n4414
g4366 and n4413 n4414_not ; n4415
g4367 nor n1021 n4415 ; n4416
g4368 nor n4415 n4416 ; n4417
g4369 nor n1021 n4416 ; n4418
g4370 nor n4417 n4418 ; n4419
g4371 nor n4316 n4319 ; n4420
g4372 nor n4333 n4420 ; n4421
g4373 nor n4308 n4313 ; n4422
g4374 and n2582_not n4307 ; n4423
g4375 nor n291 n4423 ; n4424
g4376 nor n2582 n4423 ; n4425
g4377 and n525_not n4425 ; n4426
g4378 nor n4424 n4426 ; n4427
g4379 nor n4422 n4427 ; n4428
g4380 nor n4422 n4428 ; n4429
g4381 nor n4427 n4428 ; n4430
g4382 nor n4429 n4430 ; n4431
g4383 and n2562 n2668 ; n4432
g4384 and n2578 n2776 ; n4433
g4385 and n2575_not n2666 ; n4434
g4386 nor n4433 n4434 ; n4435
g4387 and n4432_not n4435 ; n4436
g4388 and n2674_not n4436 ; n4437
g4389 and n3042_not n4436 ; n4438
g4390 nor n4437 n4438 ; n4439
g4391 and n525 n4439_not ; n4440
g4392 and n525_not n4439 ; n4441
g4393 nor n4440 n4441 ; n4442
g4394 and n4431_not n4442 ; n4443
g4395 nor n4431 n4443 ; n4444
g4396 and n4442 n4443_not ; n4445
g4397 nor n4444 n4445 ; n4446
g4398 and n2699 n3277 ; n4447
g4399 and n2566_not n2695 ; n4448
g4400 and n2554_not n2697 ; n4449
g4401 nor n4448 n4449 ; n4450
g4402 and n4447_not n4450 ; n4451
g4403 and n2690 n3332 ; n4452
g4404 and n4451 n4452_not ; n4453
g4405 nor n669 n4453 ; n4454
g4406 and n669 n4453 ; n4455
g4407 nor n4454 n4455 ; n4456
g4408 and n4446_not n4456 ; n4457
g4409 nor n4445 n4456 ; n4458
g4410 and n4444_not n4458 ; n4459
g4411 nor n4457 n4459 ; n4460
g4412 and n4421_not n4460 ; n4461
g4413 nor n4421 n4461 ; n4462
g4414 and n4460 n4461_not ; n4463
g4415 nor n4462 n4463 ; n4464
g4416 nor n4419 n4464 ; n4465
g4417 and n4419 n4463_not ; n4466
g4418 and n4462_not n4466 ; n4467
g4419 nor n4465 n4467 ; n4468
g4420 and n4408_not n4468 ; n4469
g4421 nor n4408 n4469 ; n4470
g4422 and n4468 n4469_not ; n4471
g4423 nor n4470 n4471 ; n4472
g4424 and n2560 n3750 ; n4473
g4425 and n2567 n3896 ; n4474
g4426 nor n4473 n4474 ; n4475
g4427 and n2571 n4056 ; n4476
g4428 and n4475 n4476_not ; n4477
g4429 nor n275 n4477 ; n4478
g4430 and n275 n4477 ; n4479
g4431 nor n4478 n4479 ; n4480
g4432 and n4472_not n4480 ; n4481
g4433 nor n4471 n4480 ; n4482
g4434 and n4470_not n4482 ; n4483
g4435 nor n4481 n4483 ; n4484
g4436 and n4406_not n4484 ; n4485
g4437 and n4406 n4484_not ; n4486
g4438 nor n4485 n4486 ; n4487
g4439 and n4405_not n4487 ; n4488
g4440 and n4405 n4487_not ; n4489
g4441 nor n4488 n4489 ; n4490
g4442 and n4404 n4490_not ; n4491
g4443 and n4404_not n4490 ; n4492
g4444 nor n4491 n4492 ; n4493
g4445 and n4390_not n4493 ; n4494
g4446 and n4390 n4493_not ; n4495
g4447 nor n4494 n4495 ; n4496
g4448 nor n4383 n4496 ; n4497
g4449 and n4383 n4496 ; n4498
g4450 nor n4497 n4498 ; n4499
g4451 and n4384_not n4385 ; n4500
g4452 nor n4027 n4500 ; n4501
g4453 and n4499_not n4501 ; n4502
g4454 and n4499 n4501_not ; n4503
g4455 or n4502 n4503 ; sin[5]
g4456 nor n4492 n4494 ; n4505
g4457 and n316 n1117 ; n4506
g4458 and n586 n4506 ; n4507
g4459 and n2421 n4507 ; n4508
g4460 and n2340 n4508 ; n4509
g4461 and n156 n4509 ; n4510
g4462 and n369 n4510 ; n4511
g4463 and n976 n4511 ; n4512
g4464 and n357_not n4512 ; n4513
g4465 and n253 n970 ; n4514
g4466 and n2458 n4514 ; n4515
g4467 and n3259 n4515 ; n4516
g4468 and n4513 n4516 ; n4517
g4469 and n337_not n4517 ; n4518
g4470 and n150_not n4518 ; n4519
g4471 and n172_not n4519 ; n4520
g4472 and n169_not n4520 ; n4521
g4473 and n447_not n4521 ; n4522
g4474 and n148_not n4522 ; n4523
g4475 nor n4485 n4488 ; n4524
g4476 nor n4469 n4481 ; n4525
g4477 nor n4461 n4465 ; n4526
g4478 and n2560 n3896 ; n4527
g4479 and n2571 n4054 ; n4528
g4480 nor n4527 n4528 ; n4529
g4481 and n275 n4529_not ; n4530
g4482 and n275_not n4529 ; n4531
g4483 nor n4530 n4531 ; n4532
g4484 nor n4526 n4532 ; n4533
g4485 and n4526 n4532 ; n4534
g4486 nor n4533 n4534 ; n4535
g4487 and n2802 n3750 ; n4536
g4488 and n2808 n3272 ; n4537
g4489 and n2810 n3628_not ; n4538
g4490 nor n4537 n4538 ; n4539
g4491 and n4536_not n4539 ; n4540
g4492 and n2817 n3762 ; n4541
g4493 and n4540 n4541_not ; n4542
g4494 nor n1021 n4542 ; n4543
g4495 nor n4542 n4543 ; n4544
g4496 nor n1021 n4543 ; n4545
g4497 nor n4544 n4545 ; n4546
g4498 nor n4443 n4457 ; n4547
g4499 nor n4423 n4428 ; n4548
g4500 and n2578 n4307 ; n4549
g4501 nor n291 n4549 ; n4550
g4502 and n2578 n4549_not ; n4551
g4503 and n525_not n4551 ; n4552
g4504 nor n4550 n4552 ; n4553
g4505 nor n4548 n4553 ; n4554
g4506 nor n4548 n4554 ; n4555
g4507 nor n4553 n4554 ; n4556
g4508 nor n4555 n4556 ; n4557
g4509 and n2566_not n2668 ; n4558
g4510 and n2575_not n2776 ; n4559
g4511 and n2562 n2666 ; n4560
g4512 nor n4559 n4560 ; n4561
g4513 and n4558_not n4561 ; n4562
g4514 and n2674_not n4562 ; n4563
g4515 and n3022_not n4562 ; n4564
g4516 nor n4563 n4564 ; n4565
g4517 and n525 n4565_not ; n4566
g4518 and n525_not n4565 ; n4567
g4519 nor n4566 n4567 ; n4568
g4520 and n4557_not n4568 ; n4569
g4521 nor n4557 n4569 ; n4570
g4522 and n4568 n4569_not ; n4571
g4523 nor n4570 n4571 ; n4572
g4524 and n2699 n3280_not ; n4573
g4525 and n2554_not n2695 ; n4574
g4526 and n2697 n3277 ; n4575
g4527 nor n4574 n4575 ; n4576
g4528 and n4573_not n4576 ; n4577
g4529 and n2690 n3318 ; n4578
g4530 and n4577 n4578_not ; n4579
g4531 nor n669 n4579 ; n4580
g4532 and n669 n4579 ; n4581
g4533 nor n4580 n4581 ; n4582
g4534 and n4572_not n4582 ; n4583
g4535 nor n4571 n4582 ; n4584
g4536 and n4570_not n4584 ; n4585
g4537 nor n4583 n4585 ; n4586
g4538 and n4547_not n4586 ; n4587
g4539 nor n4547 n4587 ; n4588
g4540 and n4586 n4587_not ; n4589
g4541 nor n4588 n4589 ; n4590
g4542 nor n4546 n4590 ; n4591
g4543 and n4546 n4589_not ; n4592
g4544 and n4588_not n4592 ; n4593
g4545 nor n4591 n4593 ; n4594
g4546 and n4535 n4594 ; n4595
g4547 nor n4535 n4594 ; n4596
g4548 nor n4595 n4596 ; n4597
g4549 and n4525_not n4597 ; n4598
g4550 and n4525 n4597_not ; n4599
g4551 nor n4598 n4599 ; n4600
g4552 and n4524_not n4600 ; n4601
g4553 and n4524 n4600_not ; n4602
g4554 nor n4601 n4602 ; n4603
g4555 and n4523 n4603_not ; n4604
g4556 and n4523_not n4603 ; n4605
g4557 nor n4604 n4605 ; n4606
g4558 and n4505_not n4606 ; n4607
g4559 and n4505 n4606_not ; n4608
g4560 nor n4607 n4608 ; n4609
g4561 nor n4498 n4609 ; n4610
g4562 and n4498 n4609 ; n4611
g4563 nor n4610 n4611 ; n4612
g4564 and n4499_not n4500 ; n4613
g4565 nor n4027 n4613 ; n4614
g4566 and n4612_not n4614 ; n4615
g4567 and n4612 n4614_not ; n4616
g4568 or n4615 n4616 ; sin[6]
g4569 nor n4605 n4607 ; n4618
g4570 nor n4533 n4595 ; n4619
g4571 nor n4587 n4591 ; n4620
g4572 and n2802 n3896 ; n4621
g4573 and n2808 n3628_not ; n4622
g4574 and n2810 n3750 ; n4623
g4575 nor n4622 n4623 ; n4624
g4576 and n4621_not n4624 ; n4625
g4577 and n3908_not n4625 ; n4626
g4578 and n2817_not n4625 ; n4627
g4579 nor n4626 n4627 ; n4628
g4580 and n1021 n4628_not ; n4629
g4581 and n1021_not n4628 ; n4630
g4582 nor n4629 n4630 ; n4631
g4583 and n4620_not n4631 ; n4632
g4584 and n4620 n4631_not ; n4633
g4585 nor n4632 n4633 ; n4634
g4586 nor n4569 n4583 ; n4635
g4587 nor n4549 n4554 ; n4636
g4588 and n2554_not n2668 ; n4637
g4589 and n2562 n2776 ; n4638
g4590 and n2566_not n2666 ; n4639
g4591 nor n4638 n4639 ; n4640
g4592 and n4637_not n4640 ; n4641
g4593 and n2652 n2674 ; n4642
g4594 and n4641 n4642_not ; n4643
g4595 nor n525 n4643 ; n4644
g4596 nor n4643 n4644 ; n4645
g4597 nor n525 n4644 ; n4646
g4598 nor n4645 n4646 ; n4647
g4599 nor n525 n2575 ; n4648
g4600 and n275 n291 ; n4649
g4601 nor n275 n291 ; n4650
g4602 nor n4649 n4650 ; n4651
g4603 and n4648 n4651 ; n4652
g4604 nor n4648 n4651 ; n4653
g4605 nor n4652 n4653 ; n4654
g4606 and n4647_not n4654 ; n4655
g4607 nor n4647 n4655 ; n4656
g4608 and n4654 n4655_not ; n4657
g4609 nor n4656 n4657 ; n4658
g4610 and n4636_not n4658 ; n4659
g4611 and n4636 n4658_not ; n4660
g4612 nor n4659 n4660 ; n4661
g4613 and n2699 n3272 ; n4662
g4614 and n2695 n3277 ; n4663
g4615 and n2697 n3280_not ; n4664
g4616 nor n4663 n4664 ; n4665
g4617 and n4662_not n4665 ; n4666
g4618 and n2690_not n4666 ; n4667
g4619 and n3302_not n4666 ; n4668
g4620 nor n4667 n4668 ; n4669
g4621 and n669 n4669_not ; n4670
g4622 and n669_not n4669 ; n4671
g4623 nor n4670 n4671 ; n4672
g4624 and n4661_not n4672 ; n4673
g4625 nor n4661 n4673 ; n4674
g4626 and n4672 n4673_not ; n4675
g4627 nor n4674 n4675 ; n4676
g4628 nor n4635 n4676 ; n4677
g4629 nor n4635 n4677 ; n4678
g4630 nor n4676 n4677 ; n4679
g4631 nor n4678 n4679 ; n4680
g4632 and n4634 n4680_not ; n4681
g4633 and n4634 n4681_not ; n4682
g4634 nor n4680 n4681 ; n4683
g4635 nor n4682 n4683 ; n4684
g4636 and n4619_not n4684 ; n4685
g4637 and n4619 n4684_not ; n4686
g4638 nor n4685 n4686 ; n4687
g4639 nor n4598 n4601 ; n4688
g4640 and n4687 n4688 ; n4689
g4641 nor n4687 n4688 ; n4690
g4642 nor n4689 n4690 ; n4691
g4643 and n931 n2281 ; n4692
g4644 and n4392 n4692 ; n4693
g4645 and n809 n4693 ; n4694
g4646 and n4513 n4694 ; n4695
g4647 and n129_not n4695 ; n4696
g4648 and n194_not n4696 ; n4697
g4649 and n137_not n4697 ; n4698
g4650 and n218_not n4698 ; n4699
g4651 and n1090 n4699 ; n4700
g4652 and n168_not n4700 ; n4701
g4653 and n445_not n4701 ; n4702
g4654 and n4691 n4702_not ; n4703
g4655 and n4691_not n4702 ; n4704
g4656 nor n4703 n4704 ; n4705
g4657 and n4618_not n4705 ; n4706
g4658 and n4618 n4705_not ; n4707
g4659 nor n4706 n4707 ; n4708
g4660 and n4611 n4708 ; n4709
g4661 nor n4611 n4708 ; n4710
g4662 nor n4709 n4710 ; n4711
g4663 and n4612_not n4613 ; n4712
g4664 nor n4027 n4712 ; n4713
g4665 and n4711_not n4713 ; n4714
g4666 and n4711 n4713_not ; n4715
g4667 or n4714 n4715 ; sin[7]
g4668 nor n4703 n4706 ; n4717
g4669 and n609 n2181 ; n4718
g4670 and n165 n4718 ; n4719
g4671 and n221_not n4719 ; n4720
g4672 and n219_not n4720 ; n4721
g4673 and n167_not n4721 ; n4722
g4674 and n225_not n4722 ; n4723
g4675 and n446_not n4723 ; n4724
g4676 and n111_not n4724 ; n4725
g4677 and n211_not n4725 ; n4726
g4678 and n961 n2342 ; n4727
g4679 and n979 n4727 ; n4728
g4680 and n3678 n4728 ; n4729
g4681 and n4726 n4729 ; n4730
g4682 and n408_not n4730 ; n4731
g4683 and n257_not n4731 ; n4732
g4684 and n207_not n4732 ; n4733
g4685 and n361_not n4733 ; n4734
g4686 and n224_not n4734 ; n4735
g4687 and n326_not n4735 ; n4736
g4688 and n469_not n4736 ; n4737
g4689 nor n4619 n4684 ; n4738
g4690 nor n4690 n4738 ; n4739
g4691 nor n4632 n4681 ; n4740
g4692 and n2808 n3750 ; n4741
g4693 and n2810 n3896 ; n4742
g4694 nor n4741 n4742 ; n4743
g4695 and n2817 n4056 ; n4744
g4696 and n4743 n4744_not ; n4745
g4697 nor n1021 n4745 ; n4746
g4698 nor n4745 n4746 ; n4747
g4699 nor n1021 n4746 ; n4748
g4700 nor n4747 n4748 ; n4749
g4701 nor n4673 n4677 ; n4750
g4702 nor n4636 n4658 ; n4751
g4703 nor n4655 n4751 ; n4752
g4704 and n525_not n2562 ; n4753
g4705 nor n4649 n4652 ; n4754
g4706 nor n4753 n4754 ; n4755
g4707 nor n4753 n4755 ; n4756
g4708 nor n4754 n4755 ; n4757
g4709 nor n4756 n4757 ; n4758
g4710 and n2668 n3277 ; n4759
g4711 and n2566_not n2776 ; n4760
g4712 and n2554_not n2666 ; n4761
g4713 nor n4760 n4761 ; n4762
g4714 and n4759_not n4762 ; n4763
g4715 and n2674_not n4763 ; n4764
g4716 and n3332_not n4763 ; n4765
g4717 nor n4764 n4765 ; n4766
g4718 and n525 n4766_not ; n4767
g4719 and n525_not n4766 ; n4768
g4720 nor n4767 n4768 ; n4769
g4721 and n4758_not n4769 ; n4770
g4722 and n4758 n4769_not ; n4771
g4723 nor n4770 n4771 ; n4772
g4724 and n4752_not n4772 ; n4773
g4725 nor n4752 n4773 ; n4774
g4726 and n4772 n4773_not ; n4775
g4727 nor n4774 n4775 ; n4776
g4728 and n2699 n3628_not ; n4777
g4729 and n2695 n3280_not ; n4778
g4730 and n2697 n3272 ; n4779
g4731 nor n4778 n4779 ; n4780
g4732 and n4777_not n4780 ; n4781
g4733 and n2690 n3641 ; n4782
g4734 and n4781 n4782_not ; n4783
g4735 nor n669 n4783 ; n4784
g4736 and n669 n4783 ; n4785
g4737 nor n4784 n4785 ; n4786
g4738 and n4776_not n4786 ; n4787
g4739 nor n4775 n4786 ; n4788
g4740 and n4774_not n4788 ; n4789
g4741 nor n4787 n4789 ; n4790
g4742 and n4750_not n4790 ; n4791
g4743 and n4750 n4790_not ; n4792
g4744 nor n4791 n4792 ; n4793
g4745 and n4749_not n4793 ; n4794
g4746 and n4749 n4793_not ; n4795
g4747 nor n4794 n4795 ; n4796
g4748 and n4740_not n4796 ; n4797
g4749 and n4740 n4796_not ; n4798
g4750 nor n4797 n4798 ; n4799
g4751 and n4739_not n4799 ; n4800
g4752 and n4739 n4799_not ; n4801
g4753 nor n4800 n4801 ; n4802
g4754 and n4737 n4802_not ; n4803
g4755 and n4737_not n4802 ; n4804
g4756 nor n4803 n4804 ; n4805
g4757 and n4717_not n4805 ; n4806
g4758 and n4717 n4805_not ; n4807
g4759 nor n4806 n4807 ; n4808
g4760 nor n4709 n4808 ; n4809
g4761 and n4709 n4808 ; n4810
g4762 nor n4809 n4810 ; n4811
g4763 and n4711_not n4712 ; n4812
g4764 nor n4027 n4812 ; n4813
g4765 and n4811_not n4813 ; n4814
g4766 and n4811 n4813_not ; n4815
g4767 or n4814 n4815 ; sin[8]
g4768 nor n4804 n4806 ; n4817
g4769 and n757 n809 ; n4818
g4770 and n204 n4818 ; n4819
g4771 and n3231 n4819 ; n4820
g4772 and n2432 n4820 ; n4821
g4773 and n3259 n4821 ; n4822
g4774 and n337_not n4822 ; n4823
g4775 and n327_not n4823 ; n4824
g4776 and n225_not n4824 ; n4825
g4777 and n133_not n4825 ; n4826
g4778 and n234_not n4826 ; n4827
g4779 and n356_not n4827 ; n4828
g4780 and n216_not n4828 ; n4829
g4781 nor n4791 n4794 ; n4830
g4782 nor n4755 n4770 ; n4831
g4783 and n2668 n3280_not ; n4832
g4784 and n2554_not n2776 ; n4833
g4785 and n2666 n3277 ; n4834
g4786 nor n4833 n4834 ; n4835
g4787 and n4832_not n4835 ; n4836
g4788 and n2674 n3318 ; n4837
g4789 and n4836 n4837_not ; n4838
g4790 nor n525 n4838 ; n4839
g4791 nor n4838 n4839 ; n4840
g4792 nor n525 n4839 ; n4841
g4793 nor n4840 n4841 ; n4842
g4794 and n525_not n2644 ; n4843
g4795 nor n4842 n4843 ; n4844
g4796 nor n4842 n4844 ; n4845
g4797 nor n4843 n4844 ; n4846
g4798 nor n4845 n4846 ; n4847
g4799 and n4831_not n4847 ; n4848
g4800 and n4831 n4847_not ; n4849
g4801 nor n4848 n4849 ; n4850
g4802 and n2699 n3750 ; n4851
g4803 and n2695 n3272 ; n4852
g4804 and n2697 n3628_not ; n4853
g4805 nor n4852 n4853 ; n4854
g4806 and n4851_not n4854 ; n4855
g4807 and n2690 n3762 ; n4856
g4808 and n4855 n4856_not ; n4857
g4809 nor n669 n4857 ; n4858
g4810 and n669 n4857 ; n4859
g4811 nor n4858 n4859 ; n4860
g4812 and n4850_not n4860 ; n4861
g4813 nor n4850 n4861 ; n4862
g4814 and n4860 n4861_not ; n4863
g4815 nor n4862 n4863 ; n4864
g4816 nor n4773 n4787 ; n4865
g4817 and n2808 n3896 ; n4866
g4818 and n2817 n4054 ; n4867
g4819 nor n4866 n4867 ; n4868
g4820 and n1021_not n4868 ; n4869
g4821 and n1021 n4868_not ; n4870
g4822 nor n4869 n4870 ; n4871
g4823 nor n4865 n4871 ; n4872
g4824 and n4865 n4871 ; n4873
g4825 nor n4872 n4873 ; n4874
g4826 and n4864_not n4874 ; n4875
g4827 nor n4864 n4875 ; n4876
g4828 and n4874 n4875_not ; n4877
g4829 nor n4876 n4877 ; n4878
g4830 and n4830_not n4878 ; n4879
g4831 and n4830 n4878_not ; n4880
g4832 nor n4879 n4880 ; n4881
g4833 nor n4797 n4800 ; n4882
g4834 and n4881 n4882 ; n4883
g4835 nor n4881 n4882 ; n4884
g4836 nor n4883 n4884 ; n4885
g4837 and n4829 n4885_not ; n4886
g4838 and n4829_not n4885 ; n4887
g4839 nor n4886 n4887 ; n4888
g4840 and n4817_not n4888 ; n4889
g4841 and n4817 n4888_not ; n4890
g4842 nor n4889 n4890 ; n4891
g4843 nor n4810 n4891 ; n4892
g4844 and n4810 n4891 ; n4893
g4845 nor n4892 n4893 ; n4894
g4846 and n4811_not n4812 ; n4895
g4847 nor n4027 n4895 ; n4896
g4848 and n4894_not n4896 ; n4897
g4849 and n4894 n4896_not ; n4898
g4850 or n4897 n4898 ; sin[9]
g4851 nor n4887 n4889 ; n4900
g4852 and n259 n655 ; n4901
g4853 and n476 n4901 ; n4902
g4854 and n505 n4902 ; n4903
g4855 and n210 n4903 ; n4904
g4856 and n3666 n4904 ; n4905
g4857 and n1104 n4905 ; n4906
g4858 and n3259 n4906 ; n4907
g4859 and n977 n4907 ; n4908
g4860 and n312_not n4908 ; n4909
g4861 and n192_not n4909 ; n4910
g4862 and n315_not n4910 ; n4911
g4863 nor n4830 n4878 ; n4912
g4864 nor n4884 n4912 ; n4913
g4865 nor n4872 n4875 ; n4914
g4866 nor n2566 n4753 ; n4915
g4867 and n525_not n4915 ; n4916
g4868 nor n4844 n4916 ; n4917
g4869 nor n525 n2554 ; n4918
g4870 nor n1021 n4918 ; n4919
g4871 and n1021 n4918 ; n4920
g4872 and n4753 n4920_not ; n4921
g4873 and n4919_not n4921 ; n4922
g4874 and n4753 n4922_not ; n4923
g4875 nor n4920 n4922 ; n4924
g4876 and n4919_not n4924 ; n4925
g4877 nor n4923 n4925 ; n4926
g4878 nor n4917 n4926 ; n4927
g4879 nor n4917 n4927 ; n4928
g4880 nor n4926 n4927 ; n4929
g4881 nor n4928 n4929 ; n4930
g4882 and n2668 n3272 ; n4931
g4883 and n2776 n3277 ; n4932
g4884 and n2666 n3280_not ; n4933
g4885 nor n4932 n4933 ; n4934
g4886 and n4931_not n4934 ; n4935
g4887 and n2674 n3302 ; n4936
g4888 and n4935 n4936_not ; n4937
g4889 nor n525 n4937 ; n4938
g4890 nor n525 n4938 ; n4939
g4891 nor n4937 n4938 ; n4940
g4892 nor n4939 n4940 ; n4941
g4893 nor n4930 n4941 ; n4942
g4894 nor n4930 n4942 ; n4943
g4895 nor n4941 n4942 ; n4944
g4896 nor n4943 n4944 ; n4945
g4897 nor n4831 n4847 ; n4946
g4898 nor n4861 n4946 ; n4947
g4899 and n2699 n3896 ; n4948
g4900 and n2695 n3628_not ; n4949
g4901 and n2697 n3750 ; n4950
g4902 nor n4949 n4950 ; n4951
g4903 and n4948_not n4951 ; n4952
g4904 and n2690_not n4952 ; n4953
g4905 and n3908_not n4952 ; n4954
g4906 nor n4953 n4954 ; n4955
g4907 and n669 n4955_not ; n4956
g4908 and n669_not n4955 ; n4957
g4909 nor n4956 n4957 ; n4958
g4910 and n4947_not n4958 ; n4959
g4911 nor n4947 n4959 ; n4960
g4912 and n4958 n4959_not ; n4961
g4913 nor n4960 n4961 ; n4962
g4914 nor n4945 n4962 ; n4963
g4915 and n4945 n4961_not ; n4964
g4916 and n4960_not n4964 ; n4965
g4917 nor n4963 n4965 ; n4966
g4918 and n4914_not n4966 ; n4967
g4919 and n4914 n4966_not ; n4968
g4920 nor n4967 n4968 ; n4969
g4921 and n4913_not n4969 ; n4970
g4922 and n4913 n4969_not ; n4971
g4923 nor n4970 n4971 ; n4972
g4924 and n4911 n4972_not ; n4973
g4925 and n4911_not n4972 ; n4974
g4926 nor n4973 n4974 ; n4975
g4927 and n4900_not n4975 ; n4976
g4928 and n4900 n4975_not ; n4977
g4929 nor n4976 n4977 ; n4978
g4930 nor n4893 n4978 ; n4979
g4931 and n4893 n4978 ; n4980
g4932 nor n4979 n4980 ; n4981
g4933 and n4894_not n4895 ; n4982
g4934 nor n4027 n4982 ; n4983
g4935 and n4981_not n4983 ; n4984
g4936 and n4981 n4983_not ; n4985
g4937 or n4984 n4985 ; sin[10]
g4938 nor n4974 n4976 ; n4987
g4939 and n911 n969 ; n4988
g4940 and n499 n4988 ; n4989
g4941 and n3734 n4989 ; n4990
g4942 and n636 n4990 ; n4991
g4943 and n453 n4991 ; n4992
g4944 and n336_not n4992 ; n4993
g4945 nor n4967 n4970 ; n4994
g4946 nor n4959 n4963 ; n4995
g4947 nor n4927 n4942 ; n4996
g4948 and n525_not n3277 ; n4997
g4949 and n4924_not n4997 ; n4998
g4950 and n4924 n4997_not ; n4999
g4951 nor n4998 n4999 ; n5000
g4952 and n2668 n3628_not ; n5001
g4953 and n2776 n3280_not ; n5002
g4954 and n2666 n3272 ; n5003
g4955 nor n5002 n5003 ; n5004
g4956 and n5001_not n5004 ; n5005
g4957 and n2674_not n5005 ; n5006
g4958 and n3641_not n5005 ; n5007
g4959 nor n5006 n5007 ; n5008
g4960 and n525 n5008_not ; n5009
g4961 and n525_not n5008 ; n5010
g4962 nor n5009 n5010 ; n5011
g4963 and n5000_not n5011 ; n5012
g4964 and n5000 n5011_not ; n5013
g4965 nor n5012 n5013 ; n5014
g4966 and n4996_not n5014 ; n5015
g4967 nor n4996 n5015 ; n5016
g4968 and n5014 n5015_not ; n5017
g4969 nor n5016 n5017 ; n5018
g4970 and n2695 n3750 ; n5019
g4971 and n2697 n3896 ; n5020
g4972 nor n5019 n5020 ; n5021
g4973 and n2690 n4056 ; n5022
g4974 and n5021 n5022_not ; n5023
g4975 nor n669 n5023 ; n5024
g4976 and n669 n5023 ; n5025
g4977 nor n5024 n5025 ; n5026
g4978 and n5018_not n5026 ; n5027
g4979 nor n5017 n5026 ; n5028
g4980 and n5016_not n5028 ; n5029
g4981 nor n5027 n5029 ; n5030
g4982 and n4995_not n5030 ; n5031
g4983 and n4995 n5030_not ; n5032
g4984 nor n5031 n5032 ; n5033
g4985 and n4994_not n5033 ; n5034
g4986 and n4994 n5033_not ; n5035
g4987 nor n5034 n5035 ; n5036
g4988 and n4993 n5036_not ; n5037
g4989 and n4993_not n5036 ; n5038
g4990 nor n5037 n5038 ; n5039
g4991 and n4987_not n5039 ; n5040
g4992 and n4987 n5039_not ; n5041
g4993 nor n5040 n5041 ; n5042
g4994 nor n4980 n5042 ; n5043
g4995 and n4980 n5042 ; n5044
g4996 nor n5043 n5044 ; n5045
g4997 and n4981_not n4982 ; n5046
g4998 nor n4027 n5046 ; n5047
g4999 and n5045_not n5047 ; n5048
g5000 and n5045 n5047_not ; n5049
g5001 or n5048 n5049 ; sin[11]
g5002 nor n5038 n5040 ; n5051
g5003 nor n177 n186 ; n5052
g5004 and n207_not n5052 ; n5053
g5005 and n234_not n5053 ; n5054
g5006 and n335_not n5054 ; n5055
g5007 and n2367 n5055 ; n5056
g5008 and n946 n5056 ; n5057
g5009 and n4037 n5057 ; n5058
g5010 and n2250 n5058 ; n5059
g5011 and n380 n5059 ; n5060
g5012 and n139_not n5060 ; n5061
g5013 and n134_not n5061 ; n5062
g5014 and n211_not n5062 ; n5063
g5015 nor n5031 n5034 ; n5064
g5016 nor n5015 n5027 ; n5065
g5017 and n2695 n3896 ; n5066
g5018 and n2690 n4054 ; n5067
g5019 nor n5066 n5067 ; n5068
g5020 nor n669 n5068 ; n5069
g5021 and n669 n5068 ; n5070
g5022 nor n5069 n5070 ; n5071
g5023 and n2668 n3750 ; n5072
g5024 and n2776 n3272 ; n5073
g5025 and n2666 n3628_not ; n5074
g5026 nor n5073 n5074 ; n5075
g5027 and n5072_not n5075 ; n5076
g5028 and n2674 n3762 ; n5077
g5029 and n5076 n5077_not ; n5078
g5030 nor n525 n5078 ; n5079
g5031 nor n525 n5079 ; n5080
g5032 nor n5078 n5079 ; n5081
g5033 nor n5080 n5081 ; n5082
g5034 and n5071 n5082_not ; n5083
g5035 and n5071 n5083_not ; n5084
g5036 nor n5082 n5083 ; n5085
g5037 nor n5084 n5085 ; n5086
g5038 nor n4924 n4997 ; n5087
g5039 nor n5012 n5087 ; n5088
g5040 nor n525 n3280 ; n5089
g5041 and n4997_not n5089 ; n5090
g5042 and n4997 n5089_not ; n5091
g5043 nor n5088 n5091 ; n5092
g5044 and n5090_not n5092 ; n5093
g5045 nor n5088 n5093 ; n5094
g5046 nor n5091 n5093 ; n5095
g5047 and n5090_not n5095 ; n5096
g5048 nor n5094 n5096 ; n5097
g5049 and n5086_not n5097 ; n5098
g5050 and n5086 n5097_not ; n5099
g5051 nor n5098 n5099 ; n5100
g5052 nor n5065 n5100 ; n5101
g5053 and n5065 n5100 ; n5102
g5054 nor n5101 n5102 ; n5103
g5055 and n5064_not n5103 ; n5104
g5056 and n5064 n5103_not ; n5105
g5057 nor n5104 n5105 ; n5106
g5058 and n5063 n5106_not ; n5107
g5059 and n5063_not n5106 ; n5108
g5060 nor n5107 n5108 ; n5109
g5061 and n5051_not n5109 ; n5110
g5062 and n5051 n5109_not ; n5111
g5063 nor n5110 n5111 ; n5112
g5064 nor n5044 n5112 ; n5113
g5065 and n5044 n5112 ; n5114
g5066 nor n5113 n5114 ; n5115
g5067 and n5045_not n5046 ; n5116
g5068 nor n4027 n5116 ; n5117
g5069 and n5115_not n5117 ; n5118
g5070 and n5115 n5117_not ; n5119
g5071 or n5118 n5119 ; sin[12]
g5072 nor n5108 n5110 ; n5121
g5073 nor n194 n394 ; n5122
g5074 and n255_not n5122 ; n5123
g5075 and n360_not n5123 ; n5124
g5076 and n118_not n5124 ; n5125
g5077 and n156 n5125 ; n5126
g5078 and n4002 n5126 ; n5127
g5079 and n311 n5127 ; n5128
g5080 and n2178 n5128 ; n5129
g5081 and n980 n5129 ; n5130
g5082 and n3699 n5130 ; n5131
g5083 and n196_not n5131 ; n5132
g5084 and n343_not n5132 ; n5133
g5085 and n257_not n5133 ; n5134
g5086 and n169_not n5134 ; n5135
g5087 and n142_not n5135 ; n5136
g5088 and n470_not n5136 ; n5137
g5089 and n351_not n5137 ; n5138
g5090 nor n5101 n5104 ; n5139
g5091 and n2668 n3896 ; n5140
g5092 and n2776 n3628_not ; n5141
g5093 and n2666 n3750 ; n5142
g5094 nor n5141 n5142 ; n5143
g5095 and n5140_not n5143 ; n5144
g5096 and n2674 n3908 ; n5145
g5097 and n5144 n5145_not ; n5146
g5098 nor n525 n5146 ; n5147
g5099 nor n5146 n5147 ; n5148
g5100 nor n525 n5147 ; n5149
g5101 nor n5148 n5149 ; n5150
g5102 and n669 n5089 ; n5151
g5103 nor n669 n5089 ; n5152
g5104 nor n5151 n5152 ; n5153
g5105 and n525_not n3272 ; n5154
g5106 and n5153 n5154 ; n5155
g5107 nor n5153 n5154 ; n5156
g5108 nor n5155 n5156 ; n5157
g5109 and n5150_not n5157 ; n5158
g5110 nor n5150 n5158 ; n5159
g5111 and n5157 n5158_not ; n5160
g5112 nor n5159 n5160 ; n5161
g5113 and n5095_not n5161 ; n5162
g5114 and n5095 n5161_not ; n5163
g5115 nor n5162 n5163 ; n5164
g5116 nor n5086 n5097 ; n5165
g5117 nor n5083 n5165 ; n5166
g5118 nor n5164 n5166 ; n5167
g5119 and n5164 n5166 ; n5168
g5120 nor n5167 n5168 ; n5169
g5121 and n5139_not n5169 ; n5170
g5122 and n5139 n5169_not ; n5171
g5123 nor n5170 n5171 ; n5172
g5124 and n5138_not n5172 ; n5173
g5125 and n5138 n5172_not ; n5174
g5126 nor n5121 n5174 ; n5175
g5127 and n5173_not n5175 ; n5176
g5128 nor n5121 n5176 ; n5177
g5129 nor n5173 n5176 ; n5178
g5130 and n5174_not n5178 ; n5179
g5131 nor n5177 n5179 ; n5180
g5132 and n5114_not n5180 ; n5181
g5133 and n5114 n5180_not ; n5182
g5134 nor n5181 n5182 ; n5183
g5135 and n5115_not n5116 ; n5184
g5136 nor n4027 n5184 ; n5185
g5137 and n5183_not n5185 ; n5186
g5138 and n5183 n5185_not ; n5187
g5139 or n5186 n5187 ; sin[13]
g5140 and n2367 n2433 ; n5189
g5141 and n473 n5189 ; n5190
g5142 and n967 n5190 ; n5191
g5143 and n2190 n5191 ; n5192
g5144 and n1457 n5192 ; n5193
g5145 and n983 n5193 ; n5194
g5146 and n3259 n5194 ; n5195
g5147 and n138_not n5195 ; n5196
g5148 and n176_not n5196 ; n5197
g5149 and n127_not n5197 ; n5198
g5150 and n343_not n5198 ; n5199
g5151 and n370_not n5199 ; n5200
g5152 and n336_not n5200 ; n5201
g5153 and n506_not n5201 ; n5202
g5154 nor n5167 n5170 ; n5203
g5155 nor n5095 n5161 ; n5204
g5156 nor n5158 n5204 ; n5205
g5157 nor n525 n3628 ; n5206
g5158 nor n5151 n5155 ; n5207
g5159 nor n5206 n5207 ; n5208
g5160 nor n5206 n5208 ; n5209
g5161 nor n5207 n5208 ; n5210
g5162 nor n5209 n5210 ; n5211
g5163 and n2776 n3750 ; n5212
g5164 and n2666 n3896 ; n5213
g5165 nor n5212 n5213 ; n5214
g5166 and n2674_not n5214 ; n5215
g5167 and n4056_not n5214 ; n5216
g5168 nor n5215 n5216 ; n5217
g5169 and n525 n5217_not ; n5218
g5170 and n525_not n5217 ; n5219
g5171 nor n5218 n5219 ; n5220
g5172 and n5211_not n5220 ; n5221
g5173 and n5211 n5220_not ; n5222
g5174 nor n5221 n5222 ; n5223
g5175 and n5205_not n5223 ; n5224
g5176 and n5205 n5223_not ; n5225
g5177 nor n5224 n5225 ; n5226
g5178 and n5203_not n5226 ; n5227
g5179 and n5203 n5226_not ; n5228
g5180 nor n5227 n5228 ; n5229
g5181 and n5202 n5229_not ; n5230
g5182 and n5202_not n5229 ; n5231
g5183 nor n5230 n5231 ; n5232
g5184 and n5178_not n5232 ; n5233
g5185 and n5178 n5232_not ; n5234
g5186 nor n5233 n5234 ; n5235
g5187 nor n5182 n5235 ; n5236
g5188 and n5182 n5235 ; n5237
g5189 nor n5236 n5237 ; n5238
g5190 and n5183_not n5184 ; n5239
g5191 nor n4027 n5239 ; n5240
g5192 and n5238_not n5240 ; n5241
g5193 and n5238 n5240_not ; n5242
g5194 or n5241 n5242 ; sin[14]
g5195 nor n5231 n5233 ; n5244
g5196 and n337_not n1145 ; n5245
g5197 and n328_not n5245 ; n5246
g5198 and n254_not n5246 ; n5247
g5199 and n970 n5247 ; n5248
g5200 and n344 n5248 ; n5249
g5201 and n5055 n5249 ; n5250
g5202 and n2375 n5250 ; n5251
g5203 and n1115 n5251 ; n5252
g5204 and n127_not n5252 ; n5253
g5205 and n226_not n5253 ; n5254
g5206 and n217_not n5254 ; n5255
g5207 and n356_not n5255 ; n5256
g5208 and n506_not n5256 ; n5257
g5209 and n736_not n5257 ; n5258
g5210 and n2776 n3896 ; n5259
g5211 and n2674 n4054 ; n5260
g5212 nor n5259 n5260 ; n5261
g5213 nor n525 n5261 ; n5262
g5214 nor n5261 n5262 ; n5263
g5215 nor n525 n5262 ; n5264
g5216 nor n5263 n5264 ; n5265
g5217 and n525_not n3759 ; n5266
g5218 nor n5265 n5266 ; n5267
g5219 nor n5265 n5267 ; n5268
g5220 nor n5266 n5267 ; n5269
g5221 nor n5268 n5269 ; n5270
g5222 nor n5208 n5221 ; n5271
g5223 and n5270 n5271 ; n5272
g5224 nor n5270 n5271 ; n5273
g5225 nor n5272 n5273 ; n5274
g5226 nor n5224 n5227 ; n5275
g5227 and n5274_not n5275 ; n5276
g5228 and n5274 n5275_not ; n5277
g5229 nor n5276 n5277 ; n5278
g5230 and n5258_not n5278 ; n5279
g5231 and n5258 n5278_not ; n5280
g5232 nor n5244 n5280 ; n5281
g5233 and n5279_not n5281 ; n5282
g5234 nor n5244 n5282 ; n5283
g5235 nor n5279 n5282 ; n5284
g5236 and n5280_not n5284 ; n5285
g5237 nor n5283 n5285 ; n5286
g5238 and n5237_not n5286 ; n5287
g5239 and n5237 n5286_not ; n5288
g5240 nor n5287 n5288 ; n5289
g5241 and n5238_not n5239 ; n5290
g5242 nor n4027 n5290 ; n5291
g5243 and n5289_not n5291 ; n5292
g5244 and n5289 n5291_not ; n5293
g5245 or n5292 n5293 ; sin[15]
g5246 and n638 n2313 ; n5295
g5247 and n2252 n5295 ; n5296
g5248 and n5125 n5296 ; n5297
g5249 and n233 n5297 ; n5298
g5250 and n475 n5298 ; n5299
g5251 and n3702 n5299 ; n5300
g5252 and n208_not n5300 ; n5301
g5253 and n447_not n5301 ; n5302
g5254 and n477_not n5302 ; n5303
g5255 nor n5273 n5277 ; n5304
g5256 and n3750 n5206_not ; n5305
g5257 and n525_not n5305 ; n5306
g5258 nor n5267 n5306 ; n5307
g5259 and n5304_not n5307 ; n5308
g5260 and n5304 n5307_not ; n5309
g5261 nor n5308 n5309 ; n5310
g5262 and n3896 n5206_not ; n5311
g5263 and n3896_not n5206 ; n5312
g5264 nor n5311 n5312 ; n5313
g5265 and n525_not n5313 ; n5314
g5266 and n5310 n5314_not ; n5315
g5267 and n5310_not n5314 ; n5316
g5268 nor n5315 n5316 ; n5317
g5269 nor n5303 n5317 ; n5318
g5270 and n5303 n5317 ; n5319
g5271 nor n5284 n5319 ; n5320
g5272 and n5318_not n5320 ; n5321
g5273 nor n5284 n5321 ; n5322
g5274 nor n5318 n5321 ; n5323
g5275 and n5319_not n5323 ; n5324
g5276 nor n5322 n5324 ; n5325
g5277 and n5288_not n5325 ; n5326
g5278 and n5288 n5325_not ; n5327
g5279 nor n5326 n5327 ; n5328
g5280 and n5289_not n5290 ; n5329
g5281 nor n4027 n5329 ; n5330
g5282 and n5328_not n5330 ; n5331
g5283 and n5328 n5330_not ; n5332
g5284 or n5331 n5332 ; sin[16]
g5285 and n158 n775 ; n5334
g5286 and n906 n5334 ; n5335
g5287 and n259 n5335 ; n5336
g5288 and n3243 n5336 ; n5337
g5289 and n571 n5337 ; n5338
g5290 and n980 n5338 ; n5339
g5291 and n139_not n5339 ; n5340
g5292 and n207_not n5340 ; n5341
g5293 and n297_not n5341 ; n5342
g5294 and n368_not n5342 ; n5343
g5295 and n215_not n5343 ; n5344
g5296 nor n5323 n5344 ; n5345
g5297 and n5323 n5344 ; n5346
g5298 nor n5345 n5346 ; n5347
g5299 and n5327_not n5347 ; n5348
g5300 and n5327 n5347_not ; n5349
g5301 nor n5348 n5349 ; n5350
g5302 and n5328_not n5329 ; n5351
g5303 nor n4027 n5351 ; n5352
g5304 and n5350_not n5352 ; n5353
g5305 and n5350 n5352_not ; n5354
g5306 nor n5353 n5354 ; sin[17]
g5307 and n5327 n5347 ; n5356
g5308 and n588 n2170 ; n5357
g5309 and n608 n5357 ; n5358
g5310 and n1152 n5358 ; n5359
g5311 and n1108 n5359 ; n5360
g5312 and n986 n5360 ; n5361
g5313 and n3675 n5361 ; n5362
g5314 and n176_not n5362 ; n5363
g5315 and n227_not n5363 ; n5364
g5316 and n207_not n5364 ; n5365
g5317 and n357_not n5365 ; n5366
g5318 and n238_not n5366 ; n5367
g5319 and n5345 n5367_not ; n5368
g5320 and n5345_not n5367 ; n5369
g5321 nor n5368 n5369 ; n5370
g5322 nor n5356 n5370 ; n5371
g5323 and n5356 n5369_not ; n5372
g5324 nor n5371 n5372 ; n5373
g5325 and n5350 n5351 ; n5374
g5326 nor n4027 n5374 ; n5375
g5327 and n5373_not n5375 ; n5376
g5328 and n5373 n5375_not ; n5377
g5329 or n5376 n5377 ; sin[18]
g5330 and n4392 n5247 ; n5379
g5331 and n373 n5379 ; n5380
g5332 and n2540 n5380 ; n5381
g5333 and n938 n5381 ; n5382
g5334 and n144_not n5382 ; n5383
g5335 and n152_not n5383 ; n5384
g5336 and n208_not n5384 ; n5385
g5337 and n140_not n5385 ; n5386
g5338 and n446_not n5386 ; n5387
g5339 and n298_not n5387 ; n5388
g5340 and n206_not n5388 ; n5389
g5341 and n5368_not n5389 ; n5390
g5342 and n5368 n5389_not ; n5391
g5343 nor n5390 n5391 ; n5392
g5344 nor n5372 n5392 ; n5393
g5345 and n5372 n5392 ; n5394
g5346 nor n5393 n5394 ; n5395
g5347 and n5373_not n5374 ; n5396
g5348 nor n4027 n5396 ; n5397
g5349 and n5395_not n5397 ; n5398
g5350 and n5395 n5397_not ; n5399
g5351 or n5398 n5399 ; sin[19]
g5352 and n189 n459 ; n5401
g5353 and n999 n5401 ; n5402
g5354 and n502 n5402 ; n5403
g5355 and n4726 n5403 ; n5404
g5356 and n369 n5404 ; n5405
g5357 and n194_not n5405 ; n5406
g5358 and n227_not n5406 ; n5407
g5359 and n312_not n5407 ; n5408
g5360 and n218_not n5408 ; n5409
g5361 and n213_not n5409 ; n5410
g5362 and n212_not n5410 ; n5411
g5363 and n554_not n5411 ; n5412
g5364 and n5391 n5412_not ; n5413
g5365 and n5391_not n5412 ; n5414
g5366 nor n5413 n5414 ; n5415
g5367 nor n5394 n5415 ; n5416
g5368 and n5394 n5414_not ; n5417
g5369 nor n5416 n5417 ; n5418
g5370 and n5395_not n5396 ; n5419
g5371 nor n4027 n5419 ; n5420
g5372 and n5418_not n5420 ; n5421
g5373 and n5418 n5420_not ; n5422
g5374 or n5421 n5422 ; sin[20]
g5375 and n489 n3617 ; n5424
g5376 and n444 n5424 ; n5425
g5377 and n343_not n5425 ; n5426
g5378 and n360_not n5426 ; n5427
g5379 and n5413_not n5427 ; n5428
g5380 and n5413 n5427_not ; n5429
g5381 nor n5428 n5429 ; n5430
g5382 nor n5417 n5430 ; n5431
g5383 and n5417 n5430 ; n5432
g5384 nor n5431 n5432 ; n5433
g5385 and n5418_not n5419 ; n5434
g5386 nor n4027 n5434 ; n5435
g5387 and n5433_not n5435 ; n5436
g5388 and n5433 n5435_not ; n5437
g5389 or n5436 n5437 ; sin[21]
g5390 and n444 n517 ; n5439
g5391 and n5429 n5439_not ; n5440
g5392 and n5429_not n5439 ; n5441
g5393 nor n5440 n5441 ; n5442
g5394 nor n5432 n5442 ; n5443
g5395 and n5432 n5441_not ; n5444
g5396 nor n5443 n5444 ; n5445
g5397 and n5433_not n5434 ; n5446
g5398 nor n4027 n5446 ; n5447
g5399 and n5445_not n5447 ; n5448
g5400 and n5445 n5447_not ; n5449
g5401 or n5448 n5449 ; sin[22]
g5402 and a[22]_not n71 ; n5451
g5403 nor n5440 n5444 ; n5452
g5404 and n5440 n5444 ; n5453
g5405 nor n5452 n5453 ; n5454
g5406 and n5445_not n5446 ; n5455
g5407 nor n4027 n5455 ; n5456
g5408 and n5454 n5456_not ; n5457
g5409 and n5454_not n5456 ; n5458
g5410 nor n5457 n5458 ; n5459
g5411 nand n5451_not n5459 ; sin[23]
g5412 and n5452_not n5455 ; n5461
g5413 nor n5453 n5455 ; n5462
g5414 nor n5461 n5462 ; n5463
g5415 and n5451_not n5463 ; n5464
g5416 nor n4027 n5464 ; sin[24]
g5417 not n61 ; n61_not
g5418 not n70 ; n70_not
g5419 not n53 ; n53_not
g5420 not n80 ; n80_not
g5421 not n63 ; n63_not
g5422 not n64 ; n64_not
g5423 not n91 ; n91_not
g5424 not n55 ; n55_not
g5425 not n83 ; n83_not
g5426 not n84 ; n84_not
g5427 not n93 ; n93_not
g5428 not n57 ; n57_not
g5429 not n75 ; n75_not
g5430 not n67 ; n67_not
g5431 not n86 ; n86_not
g5432 not n59 ; n59_not
g5433 not n95 ; n95_not
g5434 not n69 ; n69_not
g5435 not n97 ; n97_not
g5436 not n88 ; n88_not
g5437 not n100 ; n100_not
g5438 not n111 ; n111_not
g5439 not n300 ; n300_not
g5440 not n211 ; n211_not
g5441 not n220 ; n220_not
g5442 not n103 ; n103_not
g5443 not n140 ; n140_not
g5444 not n212 ; n212_not
g5445 not n221 ; n221_not
g5446 not n302 ; n302_not
g5447 not n213 ; n213_not
g5448 not n132 ; n132_not
g5449 not n312 ; n312_not
g5450 not n150 ; n150_not
g5451 not n114 ; n114_not
g5452 not n123 ; n123_not
g5453 not n222 ; n222_not
g5454 not n142 ; n142_not
g5455 not n214 ; n214_not
g5456 not n223 ; n223_not
g5457 not n133 ; n133_not
g5458 not n106 ; n106_not
g5459 not n313 ; n313_not
g5460 not n206 ; n206_not
g5461 not n503 ; n503_not
g5462 not n152 ; n152_not
g5463 not n224 ; n224_not
g5464 not n350 ; n350_not
g5465 not n134 ; n134_not
g5466 not n215 ; n215_not
g5467 not n324 ; n324_not
g5468 not n225 ; n225_not
g5469 not n351 ; n351_not
g5470 not n207 ; n207_not
g5471 not n315 ; n315_not
g5472 not n360 ; n360_not
g5473 not n234 ; n234_not
g5474 not n216 ; n216_not
g5475 not n504 ; n504_not
g5476 not n144 ; n144_not
g5477 not n342 ; n342_not
g5478 not n900 ; n900_not
g5479 not n405 ; n405_not
g5480 not n540 ; n540_not
g5481 not n172 ; n172_not
g5482 not n235 ; n235_not
g5483 not n127 ; n127_not
g5484 not n154 ; n154_not
g5485 not n226 ; n226_not
g5486 not n532 ; n532_not
g5487 not n361 ; n361_not
g5488 not n217 ; n217_not
g5489 not n343 ; n343_not
g5490 not n118 ; n118_not
g5491 not n415 ; n415_not
g5492 not n190 ; n190_not
g5493 not n370 ; n370_not
g5494 not n208 ; n208_not
g5495 not n271 ; n271_not
g5496 not n541 ; n541_not
g5497 not n703 ; n703_not
g5498 not n155 ; n155_not
g5499 not n254 ; n254_not
g5500 not n137 ; n137_not
g5501 not n317 ; n317_not
g5502 not n470 ; n470_not
g5503 not n146 ; n146_not
g5504 not n326 ; n326_not
g5505 not n227 ; n227_not
g5506 not n191 ; n191_not
g5507 not n335 ; n335_not
g5508 not n218 ; n218_not
g5509 not n506 ; n506_not
g5510 not n551 ; n551_not
g5511 not n722 ; n722_not
g5512 not n272 ; n272_not
g5513 not n417 ; n417_not
g5514 not n552 ; n552_not
g5515 not n129 ; n129_not
g5516 not n174 ; n174_not
g5517 not n237 ; n237_not
g5518 not n138 ; n138_not
g5519 not n228 ; n228_not
g5520 not n543 ; n543_not
g5521 not n525 ; n525_not
g5522 not n327 ; n327_not
g5523 not n192 ; n192_not
g5524 not n840 ; n840_not
g5525 not n219 ; n219_not
g5526 not n444 ; n444_not
g5527 not n291 ; n291_not
g5528 not n408 ; n408_not
g5529 not n336 ; n336_not
g5530 not n471 ; n471_not
g5531 not n255 ; n255_not
g5532 not n282 ; n282_not
g5533 not n345 ; n345_not
g5534 not n705 ; n705_not
g5535 not n832 ; n832_not
g5536 not n472 ; n472_not
g5537 not n337 ; n337_not
g5538 not n148 ; n148_not
g5539 not n445 ; n445_not
g5540 not n553 ; n553_not
g5541 not n544 ; n544_not
g5542 not n175 ; n175_not
g5543 not n670 ; n670_not
g5544 not n328 ; n328_not
g5545 not n166 ; n166_not
g5546 not n526 ; n526_not
g5547 not n139 ; n139_not
g5548 not n238 ; n238_not
g5549 not n283 ; n283_not
g5550 not n706 ; n706_not
g5551 not n715 ; n715_not
g5552 not n275 ; n275_not
g5553 not n176 ; n176_not
g5554 not n446 ; n446_not
g5555 not n554 ; n554_not
g5556 not n356 ; n356_not
g5557 not n194 ; n194_not
g5558 not n167 ; n167_not
g5559 not n257 ; n257_not
g5560 not n329 ; n329_not
g5561 not n347 ; n347_not
g5562 not n725 ; n725_not
g5563 not n833 ; n833_not
g5564 not n357 ; n357_not
g5565 not n348 ; n348_not
g5566 not n168 ; n168_not
g5567 not n258 ; n258_not
g5568 not n447 ; n447_not
g5569 not n177 ; n177_not
g5570 not n519 ; n519_not
g5571 not n186 ; n186_not
g5572 not n663 ; n663_not
g5573 not n294 ; n294_not
g5574 not n358 ; n358_not
g5575 not n367 ; n367_not
g5576 not n394 ; n394_not
g5577 not n169 ; n169_not
g5578 not n286 ; n286_not
g5579 not n736 ; n736_not
g5580 not n529 ; n529_not
g5581 not n196 ; n196_not
g5582 not n178 ; n178_not
g5583 not n277 ; n277_not
g5584 not n826 ; n826_not
g5585 not n853 ; n853_not
g5586 not n871 ; n871_not
g5587 not n188 ; n188_not
g5588 not n359 ; n359_not
g5589 not n458 ; n458_not
g5590 not n854 ; n854_not
g5591 not n494 ; n494_not
g5592 not n665 ; n665_not
g5593 not n296 ; n296_not
g5594 not n368 ; n368_not
g5595 not n692 ; n692_not
g5596 not n683 ; n683_not
g5597 not n449 ; n449_not
g5598 not n845 ; n845_not
g5599 not n548 ; n548_not
g5600 not n828 ; n828_not
g5601 not n297 ; n297_not
g5602 not n495 ; n495_not
g5603 not n468 ; n468_not
g5604 not n477 ; n477_not
g5605 not n666 ; n666_not
g5606 not n279 ; n279_not
g5607 not n891 ; n891_not
g5608 not n549 ; n549_not
g5609 not n873 ; n873_not
g5610 not n675 ; n675_not
g5611 not n864 ; n864_not
g5612 not n288 ; n288_not
g5613 not n846 ; n846_not
g5614 not n298 ; n298_not
g5615 not n469 ; n469_not
g5616 not n829 ; n829_not
g5617 not n685 ; n685_not
g5618 not n883 ; n883_not
g5619 not n865 ; n865_not
g5620 not n289 ; n289_not
g5621 not n874 ; n874_not
g5622 not n838 ; n838_not
g5623 not n677 ; n677_not
g5624 not n299 ; n299_not
g5625 not n686 ; n686_not
g5626 not n786 ; n786_not
g5627 not n669 ; n669_not
g5628 not n867 ; n867_not
g5629 not n696 ; n696_not
g5630 not n894 ; n894_not
g5631 not n885 ; n885_not
g5632 not n895 ; n895_not
g5633 not n598 ; n598_not
g5634 not n589 ; n589_not
g5635 not n697 ; n697_not
g5636 not n599 ; n599_not
g5637 not n959 ; n959_not
g5638 not n699 ; n699_not
g5639 not n897 ; n897_not
g5640 not n899 ; n899_not
g5641 not n1010 ; n1010_not
g5642 not n2000 ; n2000_not
g5643 not n2010 ; n2010_not
g5644 not n2001 ; n2001_not
g5645 not n1021 ; n1021_not
g5646 not n3001 ; n3001_not
g5647 not n2011 ; n2011_not
g5648 not n2002 ; n2002_not
g5649 not n1013 ; n1013_not
g5650 not n1130 ; n1130_not
g5651 not n1202 ; n1202_not
g5652 not n5000 ; n5000_not
g5653 not n1023 ; n1023_not
g5654 not n1041 ; n1041_not
g5655 not n3201 ; n3201_not
g5656 not n1014 ; n1014_not
g5657 not n2121 ; n2121_not
g5658 not n3102 ; n3102_not
g5659 not n1302 ; n1302_not
g5660 not n5001 ; n5001_not
g5661 not n2013 ; n2013_not
g5662 not n2022 ; n2022_not
g5663 not n1230 ; n1230_not
g5664 not n4200 ; n4200_not
g5665 not n2130 ; n2130_not
g5666 not n2031 ; n2031_not
g5667 not n4101 ; n4101_not
g5668 not n2032 ; n2032_not
g5669 not n1042 ; n1042_not
g5670 not n3022 ; n3022_not
g5671 not n3400 ; n3400_not
g5672 not n1051 ; n1051_not
g5673 not n5011 ; n5011_not
g5674 not n1501 ; n1501_not
g5675 not n2023 ; n2023_not
g5676 not n3112 ; n3112_not
g5677 not n1024 ; n1024_not
g5678 not n2122 ; n2122_not
g5679 not n1411 ; n1411_not
g5680 not n4201 ; n4201_not
g5681 not n1204 ; n1204_not
g5682 not n3500 ; n3500_not
g5683 not n2600 ; n2600_not
g5684 not n3302 ; n3302_not
g5685 not n3410 ; n3410_not
g5686 not n3212 ; n3212_not
g5687 not n3023 ; n3023_not
g5688 not n4022 ; n4022_not
g5689 not n3122 ; n3122_not
g5690 not n3320 ; n3320_not
g5691 not n3311 ; n3311_not
g5692 not n1250 ; n1250_not
g5693 not n1052 ; n1052_not
g5694 not n3401 ; n3401_not
g5695 not n1205 ; n1205_not
g5696 not n1601 ; n1601_not
g5697 not n1313 ; n1313_not
g5698 not n1007 ; n1007_not
g5699 not n4121 ; n4121_not
g5700 not n4301 ; n4301_not
g5701 not n1511 ; n1511_not
g5702 not n1520 ; n1520_not
g5703 not n1061 ; n1061_not
g5704 not n1025 ; n1025_not
g5705 not n1322 ; n1322_not
g5706 not n5030 ; n5030_not
g5707 not n1043 ; n1043_not
g5708 not n1034 ; n1034_not
g5709 not n2132 ; n2132_not
g5710 not n5022 ; n5022_not
g5711 not n1251 ; n1251_not
g5712 not n1242 ; n1242_not
g5713 not n1233 ; n1233_not
g5714 not n3042 ; n3042_not
g5715 not n1224 ; n1224_not
g5716 not n1026 ; n1026_not
g5717 not n1035 ; n1035_not
g5718 not n5103 ; n5103_not
g5719 not n1071 ; n1071_not
g5720 not n3051 ; n3051_not
g5721 not n5310 ; n5310_not
g5722 not n1341 ; n1341_not
g5723 not n3015 ; n3015_not
g5724 not n4212 ; n4212_not
g5725 not n3600 ; n3600_not
g5726 not n1512 ; n1512_not
g5727 not n1521 ; n1521_not
g5728 not n1323 ; n1323_not
g5729 not n1413 ; n1413_not
g5730 not n1431 ; n1431_not
g5731 not n1314 ; n1314_not
g5732 not n1305 ; n1305_not
g5733 not n1530 ; n1530_not
g5734 not n5202 ; n5202_not
g5735 not n5220 ; n5220_not
g5736 not n5211 ; n5211_not
g5737 not n2007 ; n2007_not
g5738 not n2124 ; n2124_not
g5739 not n2142 ; n2142_not
g5740 not n2151 ; n2151_not
g5741 not n2502 ; n2502_not
g5742 not n2025 ; n2025_not
g5743 not n2601 ; n2601_not
g5744 not n2043 ; n2043_not
g5745 not n2521 ; n2521_not
g5746 not n3016 ; n3016_not
g5747 not n1441 ; n1441_not
g5748 not n2053 ; n2053_not
g5749 not n2017 ; n2017_not
g5750 not n1702 ; n1702_not
g5751 not n1711 ; n1711_not
g5752 not n4015 ; n4015_not
g5753 not n5140 ; n5140_not
g5754 not n1810 ; n1810_not
g5755 not n1801 ; n1801_not
g5756 not n1513 ; n1513_not
g5757 not n1243 ; n1243_not
g5758 not n1009 ; n1009_not
g5759 not n2620 ; n2620_not
g5760 not n4105 ; n4105_not
g5761 not n1234 ; n1234_not
g5762 not n2611 ; n2611_not
g5763 not n2026 ; n2026_not
g5764 not n3160 ; n3160_not
g5765 not n1531 ; n1531_not
g5766 not n3106 ; n3106_not
g5767 not n3052 ; n3052_not
g5768 not n3304 ; n3304_not
g5769 not n1027 ; n1027_not
g5770 not n2530 ; n2530_not
g5771 not n3034 ; n3034_not
g5772 not n1504 ; n1504_not
g5773 not n5203 ; n5203_not
g5774 not n1621 ; n1621_not
g5775 not n4600 ; n4600_not
g5776 not n4132 ; n4132_not
g5777 not n4024 ; n4024_not
g5778 not n4501 ; n4501_not
g5779 not n5240 ; n5240_not
g5780 not n5114 ; n5114_not
g5781 not n1325 ; n1325_not
g5782 not n2108 ; n2108_not
g5783 not n4340 ; n4340_not
g5784 not n3107 ; n3107_not
g5785 not n5330 ; n5330_not
g5786 not n4322 ; n4322_not
g5787 not n1505 ; n1505_not
g5788 not n2081 ; n2081_not
g5789 not n3215 ; n3215_not
g5790 not n4241 ; n4241_not
g5791 not n3521 ; n3521_not
g5792 not n2801 ; n2801_not
g5793 not n2054 ; n2054_not
g5794 not n1721 ; n1721_not
g5795 not n1703 ; n1703_not
g5796 not n1613 ; n1613_not
g5797 not n3350 ; n3350_not
g5798 not n4421 ; n4421_not
g5799 not n3008 ; n3008_not
g5800 not n3152 ; n3152_not
g5801 not n5051 ; n5051_not
g5802 not n5420 ; n5420_not
g5803 not n3422 ; n3422_not
g5804 not n1343 ; n1343_not
g5805 not n3431 ; n3431_not
g5806 not n3035 ; n3035_not
g5807 not n2450 ; n2450_not
g5808 not n3044 ; n3044_not
g5809 not n1334 ; n1334_not
g5810 not n1352 ; n1352_not
g5811 not n1019 ; n1019_not
g5812 not n5033 ; n5033_not
g5813 not n2126 ; n2126_not
g5814 not n1370 ; n1370_not
g5815 not n2630 ; n2630_not
g5816 not n5015 ; n5015_not
g5817 not n2045 ; n2045_not
g5818 not n1442 ; n1442_not
g5819 not n5150 ; n5150_not
g5820 not n3161 ; n3161_not
g5821 not n1181 ; n1181_not
g5822 not n1082 ; n1082_not
g5823 not n2144 ; n2144_not
g5824 not n1604 ; n1604_not
g5825 not n2027 ; n2027_not
g5826 not n3332 ; n3332_not
g5827 not n4223 ; n4223_not
g5828 not n1307 ; n1307_not
g5829 not n1226 ; n1226_not
g5830 not n1316 ; n1316_not
g5831 not n2504 ; n2504_not
g5832 not n2604 ; n2604_not
g5833 not n4215 ; n4215_not
g5834 not n2136 ; n2136_not
g5835 not n1308 ; n1308_not
g5836 not n4206 ; n4206_not
g5837 not n4323 ; n4323_not
g5838 not n2640 ; n2640_not
g5839 not n4404 ; n4404_not
g5840 not n3360 ; n3360_not
g5841 not n3009 ; n3009_not
g5842 not n5304 ; n5304_not
g5843 not n1407 ; n1407_not
g5844 not n1344 ; n1344_not
g5845 not n3324 ; n3324_not
g5846 not n1353 ; n1353_not
g5847 not n1443 ; n1443_not
g5848 not n1506 ; n1506_not
g5849 not n1335 ; n1335_not
g5850 not n3603 ; n3603_not
g5851 not n3612 ; n3612_not
g5852 not n4431 ; n4431_not
g5853 not n1236 ; n1236_not
g5854 not n1263 ; n1263_not
g5855 not n5115 ; n5115_not
g5856 not n2523 ; n2523_not
g5857 not n2028 ; n2028_not
g5858 not n1803 ; n1803_not
g5859 not n1083 ; n1083_not
g5860 not n1830 ; n1830_not
g5861 not n5106 ; n5106_not
g5862 not n3216 ; n3216_not
g5863 not n4143 ; n4143_not
g5864 not n3540 ; n3540_not
g5865 not n1911 ; n1911_not
g5866 not n4260 ; n4260_not
g5867 not n1920 ; n1920_not
g5868 not n5412 ; n5412_not
g5869 not n5016 ; n5016_not
g5870 not n2622 ; n2622_not
g5871 not n4620 ; n4620_not
g5872 not n1551 ; n1551_not
g5873 not n2118 ; n2118_not
g5874 not n4233 ; n4233_not
g5875 not n1533 ; n1533_not
g5876 not n1623 ; n1623_not
g5877 not n4053 ; n4053_not
g5878 not n5232 ; n5232_not
g5879 not n3171 ; n3171_not
g5880 not n5205 ; n5205_not
g5881 not n3333 ; n3333_not
g5882 not n1272 ; n1272_not
g5883 not n5223 ; n5223_not
g5884 not n3063 ; n3063_not
g5885 not n3424 ; n3424_not
g5886 not n1354 ; n1354_not
g5887 not n3145 ; n3145_not
g5888 not n4207 ; n4207_not
g5889 not n3280 ; n3280_not
g5890 not n1336 ; n1336_not
g5891 not n4027 ; n4027_not
g5892 not n4333 ; n4333_not
g5893 not n4018 ; n4018_not
g5894 not n3505 ; n3505_not
g5895 not n5350 ; n5350_not
g5896 not n3172 ; n3172_not
g5897 not n3415 ; n3415_not
g5898 not n3370 ; n3370_not
g5899 not n3325 ; n3325_not
g5900 not n4414 ; n4414_not
g5901 not n4216 ; n4216_not
g5902 not n3550 ; n3550_not
g5903 not n1048 ; n1048_not
g5904 not n1309 ; n1309_not
g5905 not n5413 ; n5413_not
g5906 not n4432 ; n4432_not
g5907 not n1075 ; n1075_not
g5908 not n5161 ; n5161_not
g5909 not n1750 ; n1750_not
g5910 not n4090 ; n4090_not
g5911 not n1183 ; n1183_not
g5912 not n1714 ; n1714_not
g5913 not n2803 ; n2803_not
g5914 not n2632 ; n2632_not
g5915 not n4711 ; n4711_not
g5916 not n4612 ; n4612_not
g5917 not n4702 ; n4702_not
g5918 not n1615 ; n1615_not
g5919 not n1408 ; n1408_not
g5920 not n2128 ; n2128_not
g5921 not n2506 ; n2506_not
g5922 not n2164 ; n2164_not
g5923 not n4900 ; n4900_not
g5924 not n2083 ; n2083_not
g5925 not n2029 ; n2029_not
g5926 not n5008 ; n5008_not
g5927 not n5206 ; n5206_not
g5928 not n4603 ; n4603_not
g5929 not n1390 ; n1390_not
g5930 not n3028 ; n3028_not
g5931 not n4621 ; n4621_not
g5932 not n5314 ; n5314_not
g5933 not n4405 ; n4405_not
g5934 not n2156 ; n2156_not
g5935 not n5072 ; n5072_not
g5936 not n1823 ; n1823_not
g5937 not n1904 ; n1904_not
g5938 not n2660 ; n2660_not
g5939 not n4208 ; n4208_not
g5940 not n2138 ; n2138_not
g5941 not n4811 ; n4811_not
g5942 not n5090 ; n5090_not
g5943 not n4406 ; n4406_not
g5944 not n3902 ; n3902_not
g5945 not n5063 ; n5063_not
g5946 not n3344 ; n3344_not
g5947 not n2552 ; n2552_not
g5948 not n3308 ; n3308_not
g5949 not n5045 ; n5045_not
g5950 not n4802 ; n4802_not
g5951 not n3074 ; n3074_not
g5952 not n3290 ; n3290_not
g5953 not n3326 ; n3326_not
g5954 not n5441 ; n5441_not
g5955 not n1922 ; n1922_not
g5956 not n1364 ; n1364_not
g5957 not n5414 ; n5414_not
g5958 not n3461 ; n3461_not
g5959 not n3641 ; n3641_not
g5960 not n1391 ; n1391_not
g5961 not n1625 ; n1625_not
g5962 not n5018 ; n5018_not
g5963 not n5036 ; n5036_not
g5964 not n2642 ; n2642_not
g5965 not n3371 ; n3371_not
g5966 not n1409 ; n1409_not
g5967 not n1931 ; n1931_not
g5968 not n3272 ; n3272_not
g5969 not n2750 ; n2750_not
g5970 not n3209 ; n3209_not
g5971 not n1670 ; n1670_not
g5972 not n3047 ; n3047_not
g5973 not n1535 ; n1535_not
g5974 not n2831 ; n2831_not
g5975 not n1544 ; n1544_not
g5976 not n1634 ; n1634_not
g5977 not n2624 ; n2624_not
g5978 not n1382 ; n1382_not
g5979 not n4154 ; n4154_not
g5980 not n4226 ; n4226_not
g5981 not n2732 ; n2732_not
g5982 not n1175 ; n1175_not
g5983 not n1571 ; n1571_not
g5984 not n3506 ; n3506_not
g5985 not n4631 ; n4631_not
g5986 not n1553 ; n1553_not
g5987 not n5117 ; n5117_not
g5988 not n2615 ; n2615_not
g5989 not n1076 ; n1076_not
g5990 not n1805 ; n1805_not
g5991 not n4541 ; n4541_not
g5992 not n3515 ; n3515_not
g5993 not n5180 ; n5180_not
g5994 not n1751 ; n1751_not
g5995 not n1742 ; n1742_not
g5996 not n1724 ; n1724_not
g5997 not n1715 ; n1715_not
g5998 not n1328 ; n1328_not
g5999 not n1256 ; n1256_not
g6000 not n4523 ; n4523_not
g6001 not n4064 ; n4064_not
g6002 not n4028 ; n4028_not
g6003 not n4316 ; n4316_not
g6004 not n4505 ; n4505_not
g6005 not n3390 ; n3390_not
g6006 not n2571 ; n2571_not
g6007 not n3930 ; n3930_not
g6008 not n3921 ; n3921_not
g6009 not n3318 ; n3318_not
g6010 not n4128 ; n4128_not
g6011 not n3750 ; n3750_not
g6012 not n3543 ; n3543_not
g6013 not n3606 ; n3606_not
g6014 not n4191 ; n4191_not
g6015 not n2706 ; n2706_not
g6016 not n3516 ; n3516_not
g6017 not n4254 ; n4254_not
g6018 not n3471 ; n3471_not
g6019 not n4272 ; n4272_not
g6020 not n3381 ; n3381_not
g6021 not n4740 ; n4740_not
g6022 not n2607 ; n2607_not
g6023 not n2562 ; n2562_not
g6024 not n2634 ; n2634_not
g6025 not n2481 ; n2481_not
g6026 not n2508 ; n2508_not
g6027 not n4830 ; n4830_not
g6028 not n2229 ; n2229_not
g6029 not n4920 ; n4920_not
g6030 not n4911 ; n4911_not
g6031 not n2085 ; n2085_not
g6032 not n1950 ; n1950_not
g6033 not n1914 ; n1914_not
g6034 not n4470 ; n4470_not
g6035 not n4524 ; n4524_not
g6036 not n2823 ; n2823_not
g6037 not n2913 ; n2913_not
g6038 not n4614 ; n4614_not
g6039 not n2904 ; n2904_not
g6040 not n4713 ; n4713_not
g6041 not n2742 ; n2742_not
g6042 not n2751 ; n2751_not
g6043 not n2724 ; n2724_not
g6044 not n1518 ; n1518_not
g6045 not n1491 ; n1491_not
g6046 not n1356 ; n1356_not
g6047 not n5307 ; n5307_not
g6048 not n1383 ; n1383_not
g6049 not n1365 ; n1365_not
g6050 not n5325 ; n5325_not
g6051 not n1329 ; n1329_not
g6052 not n1275 ; n1275_not
g6053 not n1266 ; n1266_not
g6054 not n1257 ; n1257_not
g6055 not n5352 ; n5352_not
g6056 not n1068 ; n1068_not
g6057 not n1059 ; n1059_not
g6058 not n5433 ; n5433_not
g6059 not n5451 ; n5451_not
g6060 not n1905 ; n1905_not
g6061 not n5082 ; n5082_not
g6062 not n5064 ; n5064_not
g6063 not n5109 ; n5109_not
g6064 not n1725 ; n1725_not
g6065 not n1815 ; n1815_not
g6066 not n5145 ; n5145_not
g6067 not n1644 ; n1644_not
g6068 not n5172 ; n5172_not
g6069 not n1752 ; n1752_not
g6070 not n1716 ; n1716_not
g6071 not n4056 ; n4056_not
g6072 not n5217 ; n5217_not
g6073 not n5226 ; n5226_not
g6074 not n1635 ; n1635_not
g6075 not n1572 ; n1572_not
g6076 not n1563 ; n1563_not
g6077 not n5280 ; n5280_not
g6078 not n3066 ; n3066_not
g6079 not n3174 ; n3174_not
g6080 not n4461 ; n4461_not
g6081 not n4281 ; n4281_not
g6082 not n3084 ; n3084_not
g6083 not n4353 ; n4353_not
g6084 not n3345 ; n3345_not
g6085 not n3129 ; n3129_not
g6086 not n4362 ; n4362_not
g6087 not n4452 ; n4452_not
g6088 not n4443 ; n4443_not
g6089 not n3273 ; n3273_not
g6090 not n2815 ; n2815_not
g6091 not n2590 ; n2590_not
g6092 not n4084 ; n4084_not
g6093 not n1771 ; n1771_not
g6094 not n5173 ; n5173_not
g6095 not n2554 ; n2554_not
g6096 not n3805 ; n3805_not
g6097 not n1681 ; n1681_not
g6098 not n1960 ; n1960_not
g6099 not n1915 ; n1915_not
g6100 not n1177 ; n1177_not
g6101 not n4093 ; n4093_not
g6102 not n1942 ; n1942_not
g6103 not n1744 ; n1744_not
g6104 not n4264 ; n4264_not
g6105 not n3256 ; n3256_not
g6106 not n1951 ; n1951_not
g6107 not n5047 ; n5047_not
g6108 not n3292 ; n3292_not
g6109 not n3355 ; n3355_not
g6110 not n3490 ; n3490_not
g6111 not n5083 ; n5083_not
g6112 not n3751 ; n3751_not
g6113 not n1906 ; n1906_not
g6114 not n4336 ; n4336_not
g6115 not n1384 ; n1384_not
g6116 not n1366 ; n1366_not
g6117 not n1249 ; n1249_not
g6118 not n1186 ; n1186_not
g6119 not n3931 ; n3931_not
g6120 not n3409 ; n3409_not
g6121 not n3382 ; n3382_not
g6122 not n1258 ; n1258_not
g6123 not n1195 ; n1195_not
g6124 not n5452 ; n5452_not
g6125 not n4291 ; n4291_not
g6126 not n1690 ; n1690_not
g6127 not n3832 ; n3832_not
g6128 not n1672 ; n1672_not
g6129 not n4057 ; n4057_not
g6130 not n1627 ; n1627_not
g6131 not n1591 ; n1591_not
g6132 not n4372 ; n4372_not
g6133 not n1564 ; n1564_not
g6134 not n1537 ; n1537_not
g6135 not n3436 ; n3436_not
g6136 not n1492 ; n1492_not
g6137 not n4345 ; n4345_not
g6138 not n3643 ; n3643_not
g6139 not n2842 ; n2842_not
g6140 not n4705 ; n4705_not
g6141 not n2824 ; n2824_not
g6142 not n2806 ; n2806_not
g6143 not n2761 ; n2761_not
g6144 not n4444 ; n4444_not
g6145 not n2743 ; n2743_not
g6146 not n2734 ; n2734_not
g6147 not n4750 ; n4750_not
g6148 not n4462 ; n4462_not
g6149 not n4408 ; n4408_not
g6150 not n2932 ; n2932_not
g6151 not n3067 ; n3067_not
g6152 not n4390 ; n4390_not
g6153 not n2644 ; n2644_not
g6154 not n4570 ; n4570_not
g6155 not n4525 ; n4525_not
g6156 not n2950 ; n2950_not
g6157 not n3544 ; n3544_not
g6158 not n3562 ; n3562_not
g6159 not n4606 ; n4606_not
g6160 not n4642 ; n4642_not
g6161 not n2149 ; n2149_not
g6162 not n4147 ; n4147_not
g6163 not n3715 ; n3715_not
g6164 not n3166 ; n3166_not
g6165 not n3157 ; n3157_not
g6166 not n4831 ; n4831_not
g6167 not n3139 ; n3139_not
g6168 not n2626 ; n2626_not
g6169 not n2653 ; n2653_not
g6170 not n4813 ; n4813_not
g6171 not n2680 ; n2680_not
g6172 not n2662 ; n2662_not
g6173 not n3094 ; n3094_not
g6174 not n4085 ; n4085_not
g6175 not n4229 ; n4229_not
g6176 not n4922 ; n4922_not
g6177 not n5183 ; n5183_not
g6178 not n4931 ; n4931_not
g6179 not n4328 ; n4328_not
g6180 not n2582 ; n2582_not
g6181 not n5039 ; n5039_not
g6182 not n5327 ; n5327_not
g6183 not n4805 ; n4805_not
g6184 not n4490 ; n4490_not
g6185 not n2690 ; n2690_not
g6186 not n5345 ; n5345_not
g6187 not n4472 ; n4472_not
g6188 not n5435 ; n5435_not
g6189 not n4409 ; n4409_not
g6190 not n4319 ; n4319_not
g6191 not n4913 ; n4913_not
g6192 not n5138 ; n5138_not
g6193 not n4265 ; n4265_not
g6194 not n4832 ; n4832_not
g6195 not n5237 ; n5237_not
g6196 not n4175 ; n4175_not
g6197 not n5291 ; n5291_not
g6198 not n4148 ; n4148_not
g6199 not n4661 ; n4661_not
g6200 not n4157 ; n4157_not
g6201 not n4094 ; n4094_not
g6202 not n5174 ; n5174_not
g6203 not n4850 ; n4850_not
g6204 not n5318 ; n5318_not
g6205 not n4292 ; n4292_not
g6206 not n4463 ; n4463_not
g6207 not n4049 ; n4049_not
g6208 not n2636 ; n2636_not
g6209 not n1196 ; n1196_not
g6210 not n2960 ; n2960_not
g6211 not n2870 ; n2870_not
g6212 not n1367 ; n1367_not
g6213 not n1619 ; n1619_not
g6214 not n3635 ; n3635_not
g6215 not n1628 ; n1628_not
g6216 not n3653 ; n3653_not
g6217 not n2852 ; n2852_not
g6218 not n2843 ; n2843_not
g6219 not n1187 ; n1187_not
g6220 not n1655 ; n1655_not
g6221 not n3770 ; n3770_not
g6222 not n1178 ; n1178_not
g6223 not n2762 ; n2762_not
g6224 not n2672 ; n2672_not
g6225 not n2708 ; n2708_not
g6226 not n3392 ; n3392_not
g6227 not n3473 ; n3473_not
g6228 not n3356 ; n3356_not
g6229 not n3365 ; n3365_not
g6230 not n1358 ; n1358_not
g6231 not n3347 ; n3347_not
g6232 not n3185 ; n3185_not
g6233 not n3176 ; n3176_not
g6234 not n3095 ; n3095_not
g6235 not n3059 ; n3059_not
g6236 not n1286 ; n1286_not
g6237 not n3545 ; n3545_not
g6238 not n2942 ; n2942_not
g6239 not n1448 ; n1448_not
g6240 not n1529 ; n1529_not
g6241 not n1646 ; n1646_not
g6242 not n1790 ; n1790_not
g6243 not n1817 ; n1817_not
g6244 not n3905 ; n3905_not
g6245 not n2555 ; n2555_not
g6246 not n2528 ; n2528_not
g6247 not n1808 ; n1808_not
g6248 not n1826 ; n1826_not
g6249 not n1835 ; n1835_not
g6250 not n1862 ; n1862_not
g6251 not n2096 ; n2096_not
g6252 not n2078 ; n2078_not
g6253 not n1925 ; n1925_not
g6254 not n1970 ; n1970_not
g6255 not n1943 ; n1943_not
g6256 not n1682 ; n1682_not
g6257 not n1709 ; n1709_not
g6258 not n1736 ; n1736_not
g6259 not n2618 ; n2618_not
g6260 not n3851 ; n3851_not
g6261 not n4914 ; n4914_not
g6262 not n1863 ; n1863_not
g6263 not n1278 ; n1278_not
g6264 not n4680 ; n4680_not
g6265 not n2358 ; n2358_not
g6266 not n4446 ; n4446_not
g6267 not n1881 ; n1881_not
g6268 not n2673 ; n2673_not
g6269 not n2718 ; n2718_not
g6270 not n3078 ; n3078_not
g6271 not n2088 ; n2088_not
g6272 not n1683 ; n1683_not
g6273 not n3258 ; n3258_not
g6274 not n1962 ; n1962_not
g6275 not n3294 ; n3294_not
g6276 not n5319 ; n5319_not
g6277 not n4293 ; n4293_not
g6278 not n3339 ; n3339_not
g6279 not n1917 ; n1917_not
g6280 not n4752 ; n4752_not
g6281 not n1935 ; n1935_not
g6282 not n1944 ; n1944_not
g6283 not n2817 ; n2817_not
g6284 not n3366 ; n3366_not
g6285 not n1359 ; n1359_not
g6286 not n5328 ; n5328_not
g6287 not n1971 ; n1971_not
g6288 not n3393 ; n3393_not
g6289 not n2862 ; n2862_not
g6290 not n5238 ; n5238_not
g6291 not n1764 ; n1764_not
g6292 not n5139 ; n5139_not
g6293 not n4662 ; n4662_not
g6294 not n4851 ; n4851_not
g6295 not n2880 ; n2880_not
g6296 not n2628 ; n2628_not
g6297 not n2925 ; n2925_not
g6298 not n1809 ; n1809_not
g6299 not n1584 ; n1584_not
g6300 not n1818 ; n1818_not
g6301 not n4572 ; n4572_not
g6302 not n2646 ; n2646_not
g6303 not n5274 ; n5274_not
g6304 not n1557 ; n1557_not
g6305 not n4536 ; n4536_not
g6306 not n1746 ; n1746_not
g6307 not n1656 ; n1656_not
g6308 not n5229 ; n5229_not
g6309 not n2484 ; n2484_not
g6310 not n1647 ; n1647_not
g6311 not n5418 ; n5418_not
g6312 not n3555 ; n3555_not
g6313 not n5391 ; n5391_not
g6314 not n4257 ; n4257_not
g6315 not n3573 ; n3573_not
g6316 not n3627 ; n3627_not
g6317 not n5373 ; n5373_not
g6318 not n3870 ; n3870_not
g6319 not n4185 ; n4185_not
g6320 not n4248 ; n4248_not
g6321 not n3762 ; n3762_not
g6322 not n1296 ; n1296_not
g6323 not n3861 ; n3861_not
g6324 not n1179 ; n1179_not
g6325 not n3825 ; n3825_not
g6326 not n1269 ; n1269_not
g6327 not n4086 ; n4086_not
g6328 not n4275 ; n4275_not
g6329 not n5445 ; n5445_not
g6330 not n3456 ; n3456_not
g6331 not n5427 ; n5427_not
g6332 not n5454 ; n5454_not
g6333 not n4266 ; n4266_not
g6334 not n3942 ; n3942_not
g6335 not n2674 ; n2674_not
g6336 not n4573 ; n4573_not
g6337 not n2575 ; n2575_not
g6338 not n1666 ; n1666_not
g6339 not n2566 ; n2566_not
g6340 not n4744 ; n4744_not
g6341 not n3790 ; n3790_not
g6342 not n1657 ; n1657_not
g6343 not n3556 ; n3556_not
g6344 not n1585 ; n1585_not
g6345 not n4078 ; n4078_not
g6346 not n3628 ; n3628_not
g6347 not n5347 ; n5347_not
g6348 not n3592 ; n3592_not
g6349 not n1378 ; n1378_not
g6350 not n4636 ; n4636_not
g6351 not n4159 ; n4159_not
g6352 not n1594 ; n1594_not
g6353 not n4681 ; n4681_not
g6354 not n2836 ; n2836_not
g6355 not n4618 ; n4618_not
g6356 not n4186 ; n4186_not
g6357 not n3763 ; n3763_not
g6358 not n3916 ; n3916_not
g6359 not n2296 ; n2296_not
g6360 not n1837 ; n1837_not
g6361 not n4960 ; n4960_not
g6362 not n4924 ; n4924_not
g6363 not n5086 ; n5086_not
g6364 not n1891 ; n1891_not
g6365 not n5077 ; n5077_not
g6366 not n1873 ; n1873_not
g6367 not n1738 ; n1738_not
g6368 not n5185 ; n5185_not
g6369 not n4069 ; n4069_not
g6370 not n4717 ; n4717_not
g6371 not n2665 ; n2665_not
g6372 not n2638 ; n2638_not
g6373 not n2593 ; n2593_not
g6374 not n1765 ; n1765_not
g6375 not n1774 ; n1774_not
g6376 not n1783 ; n1783_not
g6377 not n3727 ; n3727_not
g6378 not n4861 ; n4861_not
g6379 not n3871 ; n3871_not
g6380 not n5095 ; n5095_not
g6381 not n5158 ; n5158_not
g6382 not n1297 ; n1297_not
g6383 not n4447 ; n4447_not
g6384 not n3079 ; n3079_not
g6385 not n1396 ; n1396_not
g6386 not n1189 ; n1189_not
g6387 not n4384 ; n4384_not
g6388 not n1198 ; n1198_not
g6389 not n3376 ; n3376_not
g6390 not n3394 ; n3394_not
g6391 not n3178 ; n3178_not
g6392 not n4294 ; n4294_not
g6393 not n4357 ; n4357_not
g6394 not n3358 ; n3358_not
g6395 not n4177 ; n4177_not
g6396 not n4375 ; n4375_not
g6397 not n3187 ; n3187_not
g6398 not n1369 ; n1369_not
g6399 not n3277 ; n3277_not
g6400 not n2980 ; n2980_not
g6401 not n5275 ; n5275_not
g6402 not n4817 ; n4817_not
g6403 not n3296 ; n3296_not
g6404 not n2918 ; n2918_not
g6405 not n4565 ; n4565_not
g6406 not n2909 ; n2909_not
g6407 not n3269 ; n3269_not
g6408 not n1379 ; n1379_not
g6409 not n3593 ; n3593_not
g6410 not n4178 ; n4178_not
g6411 not n3908 ; n3908_not
g6412 not n2495 ; n2495_not
g6413 not n4439 ; n4439_not
g6414 not n3836 ; n3836_not
g6415 not n4628 ; n4628_not
g6416 not n1766 ; n1766_not
g6417 not n2675 ; n2675_not
g6418 not n2693 ; n2693_not
g6419 not n4196 ; n4196_not
g6420 not n2927 ; n2927_not
g6421 not n3809 ; n3809_not
g6422 not n1928 ; n1928_not
g6423 not n3980 ; n3980_not
g6424 not n5456 ; n5456_not
g6425 not n5447 ; n5447_not
g6426 not n3953 ; n3953_not
g6427 not n4277 ; n4277_not
g6428 not n2972 ; n2972_not
g6429 not n1892 ; n1892_not
g6430 not n3377 ; n3377_not
g6431 not n5429 ; n5429_not
g6432 not n4295 ; n4295_not
g6433 not n1883 ; n1883_not
g6434 not n4547 ; n4547_not
g6435 not n1757 ; n1757_not
g6436 not n1874 ; n1874_not
g6437 not n3368 ; n3368_not
g6438 not n1865 ; n1865_not
g6439 not n1856 ; n1856_not
g6440 not n4961 ; n4961_not
g6441 not n1748 ; n1748_not
g6442 not n1586 ; n1586_not
g6443 not n1829 ; n1829_not
g6444 not n5258 ; n5258_not
g6445 not n2558 ; n2558_not
g6446 not n4637 ; n4637_not
g6447 not n4484 ; n4484_not
g6448 not n3791 ; n3791_not
g6449 not n4655 ; n4655_not
g6450 not n1289 ; n1289_not
g6451 not n3575 ; n3575_not
g6452 not n2774 ; n2774_not
g6453 not n3629 ; n3629_not
g6454 not n2783 ; n2783_not
g6455 not n2792 ; n2792_not
g6456 not n4493 ; n4493_not
g6457 not n2819 ; n2819_not
g6458 not n2873 ; n2873_not
g6459 not n3638 ; n3638_not
g6460 not n4691 ; n4691_not
g6461 not n4529 ; n4529_not
g6462 not n2756 ; n2756_not
g6463 not n3557 ; n3557_not
g6464 not n3539 ; n3539_not
g6465 not n1649 ; n1649_not
g6466 not n4619 ; n4619_not
g6467 not n4673 ; n4673_not
g6468 not n2990 ; n2990_not
g6469 not n4079 ; n4079_not
g6470 not n5375 ; n5375_not
g6471 not n4790 ; n4790_not
g6472 not n1487 ; n1487_not
g6473 not n1595 ; n1595_not
g6474 not n1676 ; n1676_not
g6475 not n2586 ; n2586_not
g6476 not n5097 ; n5097_not
g6477 not n1695 ; n1695_not
g6478 not n4782 ; n4782_not
g6479 not n5439 ; n5439_not
g6480 not n2649 ; n2649_not
g6481 not n1857 ; n1857_not
g6482 not n1578 ; n1578_not
g6483 not n3747 ; n3747_not
g6484 not n5286 ; n5286_not
g6485 not n3387 ; n3387_not
g6486 not n4296 ; n4296_not
g6487 not n1929 ; n1929_not
g6488 not n3945 ; n3945_not
g6489 not n1983 ; n1983_not
g6490 not n3585 ; n3585_not
g6491 not n1992 ; n1992_not
g6492 not n4737 ; n4737_not
g6493 not n5178 ; n5178_not
g6494 not n3756 ; n3756_not
g6495 not n3909 ; n3909_not
g6496 not n2757 ; n2757_not
g6497 not n2739 ; n2739_not
g6498 not n4773 ; n4773_not
g6499 not n4386 ; n4386_not
g6500 not n3288 ; n3288_not
g6501 not n3783 ; n3783_not
g6502 not n1659 ; n1659_not
g6503 not n4647 ; n4647_not
g6504 not n3576 ; n3576_not
g6505 not n3864 ; n3864_not
g6506 not n5169 ; n5169_not
g6507 not n4476 ; n4476_not
g6508 not n5367 ; n5367_not
g6509 not n1668 ; n1668_not
g6510 not n2955 ; n2955_not
g6511 not n1758 ; n1758_not
g6512 not n4197 ; n4197_not
g6513 not n3936 ; n3936_not
g6514 not n4557 ; n4557_not
g6515 not n2856 ; n2856_not
g6516 not n1389 ; n1389_not
g6517 not n1398 ; n1398_not
g6518 not n1759 ; n1759_not
g6519 not n5368 ; n5368_not
g6520 not n5089 ; n5089_not
g6521 not n5278 ; n5278_not
g6522 not n5395 ; n5395_not
g6523 not n1597 ; n1597_not
g6524 not n1579 ; n1579_not
g6525 not n1399 ; n1399_not
g6526 not n4981 ; n4981_not
g6527 not n1786 ; n1786_not
g6528 not n2929 ; n2929_not
g6529 not n4972 ; n4972_not
g6530 not n4549 ; n4549_not
g6531 not n4558 ; n4558_not
g6532 not n3937 ; n3937_not
g6533 not n2965 ; n2965_not
g6534 not n2839 ; n2839_not
g6535 not n2893 ; n2893_not
g6536 not n4936 ; n4936_not
g6537 not n2857 ; n2857_not
g6538 not n4684 ; n4684_not
g6539 not n4774 ; n4774_not
g6540 not n4864 ; n4864_not
g6541 not n2686 ; n2686_not
g6542 not n2578 ; n2578_not
g6543 not n4837 ; n4837_not
g6544 not n2596 ; n2596_not
g6545 not n1984 ; n1984_not
g6546 not n3379 ; n3379_not
g6547 not n3388 ; n3388_not
g6548 not n4369 ; n4369_not
g6549 not n4378 ; n4378_not
g6550 not n3496 ; n3496_not
g6551 not n3946 ; n3946_not
g6552 not n3784 ; n3784_not
g6553 not n3199 ; n3199_not
g6554 not n3973 ; n3973_not
g6555 not n3568 ; n3568_not
g6556 not n3586 ; n3586_not
g6557 not n1993 ; n1993_not
g6558 not n3649 ; n3649_not
g6559 not n3775 ; n3775_not
g6560 not n4739 ; n4739_not
g6561 not n2696 ; n2696_not
g6562 not n4793 ; n4793_not
g6563 not n3488 ; n3488_not
g6564 not n1688 ; n1688_not
g6565 not n4766 ; n4766_not
g6566 not n2759 ; n2759_not
g6567 not n2849 ; n2849_not
g6568 not n2867 ; n2867_not
g6569 not n4658 ; n4658_not
g6570 not n5288 ; n5288_not
g6571 not n3299 ; n3299_not
g6572 not n5279 ; n5279_not
g6573 not n3794 ; n3794_not
g6574 not n2939 ; n2939_not
g6575 not n4487 ; n4487_not
g6576 not n5369 ; n5369_not
g6577 not n4469 ; n4469_not
g6578 not n4955 ; n4955_not
g6579 not n4919 ; n4919_not
g6580 not n4829 ; n4829_not
g6581 not n3875 ; n3875_not
g6582 not n3938 ; n3938_not
g6583 not n1976 ; n1976_not
g6584 not n1787 ; n1787_not
g6585 not n3893 ; n3893_not
g6586 not n2597 ; n2597_not
g6587 not n4847 ; n4847_not
g6588 not n4856 ; n4856_not
g6589 not n4587 ; n4587_not
g6590 not n4578 ; n4578_not
g6591 not n3759 ; n3759_not
g6592 not n4947 ; n4947_not
g6593 not n4569 ; n4569_not
g6594 not n3876 ; n3876_not
g6595 not n1797 ; n1797_not
g6596 not n3498 ; n3498_not
g6597 not n1869 ; n1869_not
g6598 not n5289 ; n5289_not
g6599 not n1878 ; n1878_not
g6600 not n4983 ; n4983_not
g6601 not n1977 ; n1977_not
g6602 not n2895 ; n2895_not
g6603 not n1995 ; n1995_not
g6604 not n3984 ; n3984_not
g6605 not n1986 ; n1986_not
g6606 not n3399 ; n3399_not
g6607 not n3957 ; n3957_not
g6608 not n4776 ; n4776_not
g6609 not n1698 ; n1698_not
g6610 not n4749 ; n4749_not
g6611 not n1599 ; n1599_not
g6612 not n1689 ; n1689_not
g6613 not n4875 ; n4875_not
g6614 not n5397 ; n5397_not
g6615 not n4758 ; n4758_not
g6616 not n2769 ; n2769_not
g6617 not n4885 ; n4885_not
g6618 not n4777 ; n4777_not
g6619 not n4894 ; n4894_not
g6620 not n4975 ; n4975_not
g6621 not n1879 ; n1879_not
g6622 not n4759 ; n4759_not
g6623 not n3499 ; n3499_not
g6624 not n5389 ; n5389_not
g6625 not n1978 ; n1978_not
g6626 not n4966 ; n4966_not
g6627 not n4669 ; n4669_not
g6628 not n4948 ; n4948_not
g6629 not n3589 ; n3589_not
g6630 not n4588 ; n4588_not
g6631 not n4597 ; n4597_not
g6632 not n4993 ; n4993_not
g6633 not n2689 ; n2689_not
g6634 not n4868 ; n4868_not
g6635 not n4796 ; n4796_not
g6636 not n4994 ; n4994_not
g6637 not n1898 ; n1898_not
g6638 not n1997 ; n1997_not
g6639 not n3896 ; n3896_not
g6640 not n4769 ; n4769_not
g6641 not n1799 ; n1799_not
g6642 not n4499 ; n4499_not
g6643 not n1889 ; n1889_not
g6644 not n2798 ; n2798_not
g6645 not n2888 ; n2888_not
g6646 not n4589 ; n4589_not
g6647 not n2897 ; n2897_not
g6648 not n3789 ; n3789_not
g6649 not n3798 ; n3798_not
g6650 not n3897 ; n3897_not
g6651 not a[0] ; a[0]_not
g6652 not n4995 ; n4995_not
g6653 not n1989 ; n1989_not
g6654 not n1899 ; n1899_not
g6655 not n4959 ; n4959_not
g6656 not n2997 ; n2997_not
g6657 not n4896 ; n4896_not
g6658 not n4878 ; n4878_not
g6659 not n2979 ; n2979_not
g6660 not n4987 ; n4987_not
g6661 not n4996 ; n4996_not
g6662 not n2989 ; n2989_not
g6663 not n4969 ; n4969_not
g6664 not n4888 ; n4888_not
g6665 not a[1] ; a[1]_not
g6666 not n4997 ; n4997_not
g6667 not n4799 ; n4799_not
g6668 not a[3] ; a[3]_not
g6669 not n3999 ; n3999_not
g6670 not a[4] ; a[4]_not
g6671 not a[5] ; a[5]_not
g6672 not a[6] ; a[6]_not
g6673 not a[7] ; a[7]_not
g6674 not a[8] ; a[8]_not
g6675 not a[9] ; a[9]_not
g6676 not a[10] ; a[10]_not
g6677 not a[20] ; a[20]_not
g6678 not a[11] ; a[11]_not
g6679 not a[12] ; a[12]_not
g6680 not a[21] ; a[21]_not
g6681 not a[13] ; a[13]_not
g6682 not a[22] ; a[22]_not
g6683 not a[23] ; a[23]_not
g6684 not a[14] ; a[14]_not
g6685 not a[15] ; a[15]_not
g6686 not a[16] ; a[16]_not
g6687 not a[17] ; a[17]_not
g6688 not a[18] ; a[18]_not
g6689 not a[19] ; a[19]_not
