name dec
i count[0]
i count[1]
i count[2]
i count[3]
i count[4]
i count[5]
i count[6]
i count[7]

g1 and count[4]_not count[5]_not ; n265
g2 and count[6]_not count[7] ; n266
g3 and n265 n266 ; n267
g4 and count[0]_not count[2]_not ; n268
g5 and count[1]_not count[3]_not ; n269
g6 and n268 n269 ; n270
g7 and n267 n270 ; selectp1[0]
g8 and count[0] count[2]_not ; n272
g9 and n269 n272 ; n273
g10 and n267 n273 ; selectp1[1]
g11 and count[1] count[3]_not ; n275
g12 and n268 n275 ; n276
g13 and n267 n276 ; selectp1[2]
g14 and n272 n275 ; n278
g15 and n267 n278 ; selectp1[3]
g16 and count[0]_not count[2] ; n280
g17 and n269 n280 ; n281
g18 and n267 n281 ; selectp1[4]
g19 and count[0] count[2] ; n283
g20 and n269 n283 ; n284
g21 and n267 n284 ; selectp1[5]
g22 and n275 n280 ; n286
g23 and n267 n286 ; selectp1[6]
g24 and n275 n283 ; n288
g25 and n267 n288 ; selectp1[7]
g26 and count[1]_not count[3] ; n290
g27 and n268 n290 ; n291
g28 and n267 n291 ; selectp1[8]
g29 and n272 n290 ; n293
g30 and n267 n293 ; selectp1[9]
g31 and count[1] count[3] ; n295
g32 and n268 n295 ; n296
g33 and n267 n296 ; selectp1[10]
g34 and n272 n295 ; n298
g35 and n267 n298 ; selectp1[11]
g36 and n280 n290 ; n300
g37 and n267 n300 ; selectp1[12]
g38 and n283 n290 ; n302
g39 and n267 n302 ; selectp1[13]
g40 and n280 n295 ; n304
g41 and n267 n304 ; selectp1[14]
g42 and n283 n295 ; n306
g43 and n267 n306 ; selectp1[15]
g44 and count[4] count[5]_not ; n308
g45 and n266 n308 ; n309
g46 and n270 n309 ; selectp1[16]
g47 and n273 n309 ; selectp1[17]
g48 and n276 n309 ; selectp1[18]
g49 and n278 n309 ; selectp1[19]
g50 and n281 n309 ; selectp1[20]
g51 and n284 n309 ; selectp1[21]
g52 and n286 n309 ; selectp1[22]
g53 and n288 n309 ; selectp1[23]
g54 and n291 n309 ; selectp1[24]
g55 and n293 n309 ; selectp1[25]
g56 and n296 n309 ; selectp1[26]
g57 and n298 n309 ; selectp1[27]
g58 and n300 n309 ; selectp1[28]
g59 and n302 n309 ; selectp1[29]
g60 and n304 n309 ; selectp1[30]
g61 and n306 n309 ; selectp1[31]
g62 and count[4]_not count[5] ; n326
g63 and n266 n326 ; n327
g64 and n270 n327 ; selectp1[32]
g65 and n273 n327 ; selectp1[33]
g66 and n276 n327 ; selectp1[34]
g67 and n278 n327 ; selectp1[35]
g68 and n281 n327 ; selectp1[36]
g69 and n284 n327 ; selectp1[37]
g70 and n286 n327 ; selectp1[38]
g71 and n288 n327 ; selectp1[39]
g72 and n291 n327 ; selectp1[40]
g73 and n293 n327 ; selectp1[41]
g74 and n296 n327 ; selectp1[42]
g75 and n298 n327 ; selectp1[43]
g76 and n300 n327 ; selectp1[44]
g77 and n302 n327 ; selectp1[45]
g78 and n304 n327 ; selectp1[46]
g79 and n306 n327 ; selectp1[47]
g80 and count[4] count[5] ; n344
g81 and n266 n344 ; n345
g82 and n270 n345 ; selectp1[48]
g83 and n273 n345 ; selectp1[49]
g84 and n276 n345 ; selectp1[50]
g85 and n278 n345 ; selectp1[51]
g86 and n281 n345 ; selectp1[52]
g87 and n284 n345 ; selectp1[53]
g88 and n286 n345 ; selectp1[54]
g89 and n288 n345 ; selectp1[55]
g90 and n291 n345 ; selectp1[56]
g91 and n293 n345 ; selectp1[57]
g92 and n296 n345 ; selectp1[58]
g93 and n298 n345 ; selectp1[59]
g94 and n300 n345 ; selectp1[60]
g95 and n302 n345 ; selectp1[61]
g96 and n304 n345 ; selectp1[62]
g97 and n306 n345 ; selectp1[63]
g98 and count[6] count[7] ; n362
g99 and n265 n362 ; n363
g100 and n270 n363 ; selectp1[64]
g101 and n273 n363 ; selectp1[65]
g102 and n276 n363 ; selectp1[66]
g103 and n278 n363 ; selectp1[67]
g104 and n281 n363 ; selectp1[68]
g105 and n284 n363 ; selectp1[69]
g106 and n286 n363 ; selectp1[70]
g107 and n288 n363 ; selectp1[71]
g108 and n291 n363 ; selectp1[72]
g109 and n293 n363 ; selectp1[73]
g110 and n296 n363 ; selectp1[74]
g111 and n298 n363 ; selectp1[75]
g112 and n300 n363 ; selectp1[76]
g113 and n302 n363 ; selectp1[77]
g114 and n304 n363 ; selectp1[78]
g115 and n306 n363 ; selectp1[79]
g116 and n308 n362 ; n380
g117 and n270 n380 ; selectp1[80]
g118 and n273 n380 ; selectp1[81]
g119 and n276 n380 ; selectp1[82]
g120 and n278 n380 ; selectp1[83]
g121 and n281 n380 ; selectp1[84]
g122 and n284 n380 ; selectp1[85]
g123 and n286 n380 ; selectp1[86]
g124 and n288 n380 ; selectp1[87]
g125 and n291 n380 ; selectp1[88]
g126 and n293 n380 ; selectp1[89]
g127 and n296 n380 ; selectp1[90]
g128 and n298 n380 ; selectp1[91]
g129 and n300 n380 ; selectp1[92]
g130 and n302 n380 ; selectp1[93]
g131 and n304 n380 ; selectp1[94]
g132 and n306 n380 ; selectp1[95]
g133 and n326 n362 ; n397
g134 and n270 n397 ; selectp1[96]
g135 and n273 n397 ; selectp1[97]
g136 and n276 n397 ; selectp1[98]
g137 and n278 n397 ; selectp1[99]
g138 and n281 n397 ; selectp1[100]
g139 and n284 n397 ; selectp1[101]
g140 and n286 n397 ; selectp1[102]
g141 and n288 n397 ; selectp1[103]
g142 and n291 n397 ; selectp1[104]
g143 and n293 n397 ; selectp1[105]
g144 and n296 n397 ; selectp1[106]
g145 and n298 n397 ; selectp1[107]
g146 and n300 n397 ; selectp1[108]
g147 and n302 n397 ; selectp1[109]
g148 and n304 n397 ; selectp1[110]
g149 and n306 n397 ; selectp1[111]
g150 and n344 n362 ; n414
g151 and n270 n414 ; selectp1[112]
g152 and n273 n414 ; selectp1[113]
g153 and n276 n414 ; selectp1[114]
g154 and n278 n414 ; selectp1[115]
g155 and n281 n414 ; selectp1[116]
g156 and n284 n414 ; selectp1[117]
g157 and n286 n414 ; selectp1[118]
g158 and n288 n414 ; selectp1[119]
g159 and n291 n414 ; selectp1[120]
g160 and n293 n414 ; selectp1[121]
g161 and n296 n414 ; selectp1[122]
g162 and n298 n414 ; selectp1[123]
g163 and n300 n414 ; selectp1[124]
g164 and n302 n414 ; selectp1[125]
g165 and n304 n414 ; selectp1[126]
g166 and n306 n414 ; selectp1[127]
g167 and count[6]_not count[7]_not ; n431
g168 and n265 n431 ; n432
g169 and n270 n432 ; selectp2[0]
g170 and n273 n432 ; selectp2[1]
g171 and n276 n432 ; selectp2[2]
g172 and n278 n432 ; selectp2[3]
g173 and n281 n432 ; selectp2[4]
g174 and n284 n432 ; selectp2[5]
g175 and n286 n432 ; selectp2[6]
g176 and n288 n432 ; selectp2[7]
g177 and n291 n432 ; selectp2[8]
g178 and n293 n432 ; selectp2[9]
g179 and n296 n432 ; selectp2[10]
g180 and n298 n432 ; selectp2[11]
g181 and n300 n432 ; selectp2[12]
g182 and n302 n432 ; selectp2[13]
g183 and n304 n432 ; selectp2[14]
g184 and n306 n432 ; selectp2[15]
g185 and n308 n431 ; n449
g186 and n270 n449 ; selectp2[16]
g187 and n273 n449 ; selectp2[17]
g188 and n276 n449 ; selectp2[18]
g189 and n278 n449 ; selectp2[19]
g190 and n281 n449 ; selectp2[20]
g191 and n284 n449 ; selectp2[21]
g192 and n286 n449 ; selectp2[22]
g193 and n288 n449 ; selectp2[23]
g194 and n291 n449 ; selectp2[24]
g195 and n293 n449 ; selectp2[25]
g196 and n296 n449 ; selectp2[26]
g197 and n298 n449 ; selectp2[27]
g198 and n300 n449 ; selectp2[28]
g199 and n302 n449 ; selectp2[29]
g200 and n304 n449 ; selectp2[30]
g201 and n306 n449 ; selectp2[31]
g202 and n326 n431 ; n466
g203 and n270 n466 ; selectp2[32]
g204 and n273 n466 ; selectp2[33]
g205 and n276 n466 ; selectp2[34]
g206 and n278 n466 ; selectp2[35]
g207 and n281 n466 ; selectp2[36]
g208 and n284 n466 ; selectp2[37]
g209 and n286 n466 ; selectp2[38]
g210 and n288 n466 ; selectp2[39]
g211 and n291 n466 ; selectp2[40]
g212 and n293 n466 ; selectp2[41]
g213 and n296 n466 ; selectp2[42]
g214 and n298 n466 ; selectp2[43]
g215 and n300 n466 ; selectp2[44]
g216 and n302 n466 ; selectp2[45]
g217 and n304 n466 ; selectp2[46]
g218 and n306 n466 ; selectp2[47]
g219 and n344 n431 ; n483
g220 and n270 n483 ; selectp2[48]
g221 and n273 n483 ; selectp2[49]
g222 and n276 n483 ; selectp2[50]
g223 and n278 n483 ; selectp2[51]
g224 and n281 n483 ; selectp2[52]
g225 and n284 n483 ; selectp2[53]
g226 and n286 n483 ; selectp2[54]
g227 and n288 n483 ; selectp2[55]
g228 and n291 n483 ; selectp2[56]
g229 and n293 n483 ; selectp2[57]
g230 and n296 n483 ; selectp2[58]
g231 and n298 n483 ; selectp2[59]
g232 and n300 n483 ; selectp2[60]
g233 and n302 n483 ; selectp2[61]
g234 and n304 n483 ; selectp2[62]
g235 and n306 n483 ; selectp2[63]
g236 and count[6] count[7]_not ; n500
g237 and n265 n500 ; n501
g238 and n270 n501 ; selectp2[64]
g239 and n273 n501 ; selectp2[65]
g240 and n276 n501 ; selectp2[66]
g241 and n278 n501 ; selectp2[67]
g242 and n281 n501 ; selectp2[68]
g243 and n284 n501 ; selectp2[69]
g244 and n286 n501 ; selectp2[70]
g245 and n288 n501 ; selectp2[71]
g246 and n291 n501 ; selectp2[72]
g247 and n293 n501 ; selectp2[73]
g248 and n296 n501 ; selectp2[74]
g249 and n298 n501 ; selectp2[75]
g250 and n300 n501 ; selectp2[76]
g251 and n302 n501 ; selectp2[77]
g252 and n304 n501 ; selectp2[78]
g253 and n306 n501 ; selectp2[79]
g254 and n308 n500 ; n518
g255 and n270 n518 ; selectp2[80]
g256 and n273 n518 ; selectp2[81]
g257 and n276 n518 ; selectp2[82]
g258 and n278 n518 ; selectp2[83]
g259 and n281 n518 ; selectp2[84]
g260 and n284 n518 ; selectp2[85]
g261 and n286 n518 ; selectp2[86]
g262 and n288 n518 ; selectp2[87]
g263 and n291 n518 ; selectp2[88]
g264 and n293 n518 ; selectp2[89]
g265 and n296 n518 ; selectp2[90]
g266 and n298 n518 ; selectp2[91]
g267 and n300 n518 ; selectp2[92]
g268 and n302 n518 ; selectp2[93]
g269 and n304 n518 ; selectp2[94]
g270 and n306 n518 ; selectp2[95]
g271 and n326 n500 ; n535
g272 and n270 n535 ; selectp2[96]
g273 and n273 n535 ; selectp2[97]
g274 and n276 n535 ; selectp2[98]
g275 and n278 n535 ; selectp2[99]
g276 and n281 n535 ; selectp2[100]
g277 and n284 n535 ; selectp2[101]
g278 and n286 n535 ; selectp2[102]
g279 and n288 n535 ; selectp2[103]
g280 and n291 n535 ; selectp2[104]
g281 and n293 n535 ; selectp2[105]
g282 and n296 n535 ; selectp2[106]
g283 and n298 n535 ; selectp2[107]
g284 and n300 n535 ; selectp2[108]
g285 and n302 n535 ; selectp2[109]
g286 and n304 n535 ; selectp2[110]
g287 and n306 n535 ; selectp2[111]
g288 and n344 n500 ; n552
g289 and n270 n552 ; selectp2[112]
g290 and n273 n552 ; selectp2[113]
g291 and n276 n552 ; selectp2[114]
g292 and n278 n552 ; selectp2[115]
g293 and n281 n552 ; selectp2[116]
g294 and n284 n552 ; selectp2[117]
g295 and n286 n552 ; selectp2[118]
g296 and n288 n552 ; selectp2[119]
g297 and n291 n552 ; selectp2[120]
g298 and n293 n552 ; selectp2[121]
g299 and n296 n552 ; selectp2[122]
g300 and n298 n552 ; selectp2[123]
g301 and n300 n552 ; selectp2[124]
g302 and n302 n552 ; selectp2[125]
g303 and n304 n552 ; selectp2[126]
g304 and n306 n552 ; selectp2[127]
g305 not count[4] ; count[4]_not
g306 not count[5] ; count[5]_not
g307 not count[6] ; count[6]_not
g308 not count[0] ; count[0]_not
g309 not count[2] ; count[2]_not
g310 not count[1] ; count[1]_not
g311 not count[3] ; count[3]_not
g312 not count[7] ; count[7]_not
o selectp1[0]
o selectp1[1]
o selectp1[2]
o selectp1[3]
o selectp1[4]
o selectp1[5]
o selectp1[6]
o selectp1[7]
o selectp1[8]
o selectp1[9]
o selectp1[10]
o selectp1[11]
o selectp1[12]
o selectp1[13]
o selectp1[14]
o selectp1[15]
o selectp1[16]
o selectp1[17]
o selectp1[18]
o selectp1[19]
o selectp1[20]
o selectp1[21]
o selectp1[22]
o selectp1[23]
o selectp1[24]
o selectp1[25]
o selectp1[26]
o selectp1[27]
o selectp1[28]
o selectp1[29]
o selectp1[30]
o selectp1[31]
o selectp1[32]
o selectp1[33]
o selectp1[34]
o selectp1[35]
o selectp1[36]
o selectp1[37]
o selectp1[38]
o selectp1[39]
o selectp1[40]
o selectp1[41]
o selectp1[42]
o selectp1[43]
o selectp1[44]
o selectp1[45]
o selectp1[46]
o selectp1[47]
o selectp1[48]
o selectp1[49]
o selectp1[50]
o selectp1[51]
o selectp1[52]
o selectp1[53]
o selectp1[54]
o selectp1[55]
o selectp1[56]
o selectp1[57]
o selectp1[58]
o selectp1[59]
o selectp1[60]
o selectp1[61]
o selectp1[62]
o selectp1[63]
o selectp1[64]
o selectp1[65]
o selectp1[66]
o selectp1[67]
o selectp1[68]
o selectp1[69]
o selectp1[70]
o selectp1[71]
o selectp1[72]
o selectp1[73]
o selectp1[74]
o selectp1[75]
o selectp1[76]
o selectp1[77]
o selectp1[78]
o selectp1[79]
o selectp1[80]
o selectp1[81]
o selectp1[82]
o selectp1[83]
o selectp1[84]
o selectp1[85]
o selectp1[86]
o selectp1[87]
o selectp1[88]
o selectp1[89]
o selectp1[90]
o selectp1[91]
o selectp1[92]
o selectp1[93]
o selectp1[94]
o selectp1[95]
o selectp1[96]
o selectp1[97]
o selectp1[98]
o selectp1[99]
o selectp1[100]
o selectp1[101]
o selectp1[102]
o selectp1[103]
o selectp1[104]
o selectp1[105]
o selectp1[106]
o selectp1[107]
o selectp1[108]
o selectp1[109]
o selectp1[110]
o selectp1[111]
o selectp1[112]
o selectp1[113]
o selectp1[114]
o selectp1[115]
o selectp1[116]
o selectp1[117]
o selectp1[118]
o selectp1[119]
o selectp1[120]
o selectp1[121]
o selectp1[122]
o selectp1[123]
o selectp1[124]
o selectp1[125]
o selectp1[126]
o selectp1[127]
o selectp2[0]
o selectp2[1]
o selectp2[2]
o selectp2[3]
o selectp2[4]
o selectp2[5]
o selectp2[6]
o selectp2[7]
o selectp2[8]
o selectp2[9]
o selectp2[10]
o selectp2[11]
o selectp2[12]
o selectp2[13]
o selectp2[14]
o selectp2[15]
o selectp2[16]
o selectp2[17]
o selectp2[18]
o selectp2[19]
o selectp2[20]
o selectp2[21]
o selectp2[22]
o selectp2[23]
o selectp2[24]
o selectp2[25]
o selectp2[26]
o selectp2[27]
o selectp2[28]
o selectp2[29]
o selectp2[30]
o selectp2[31]
o selectp2[32]
o selectp2[33]
o selectp2[34]
o selectp2[35]
o selectp2[36]
o selectp2[37]
o selectp2[38]
o selectp2[39]
o selectp2[40]
o selectp2[41]
o selectp2[42]
o selectp2[43]
o selectp2[44]
o selectp2[45]
o selectp2[46]
o selectp2[47]
o selectp2[48]
o selectp2[49]
o selectp2[50]
o selectp2[51]
o selectp2[52]
o selectp2[53]
o selectp2[54]
o selectp2[55]
o selectp2[56]
o selectp2[57]
o selectp2[58]
o selectp2[59]
o selectp2[60]
o selectp2[61]
o selectp2[62]
o selectp2[63]
o selectp2[64]
o selectp2[65]
o selectp2[66]
o selectp2[67]
o selectp2[68]
o selectp2[69]
o selectp2[70]
o selectp2[71]
o selectp2[72]
o selectp2[73]
o selectp2[74]
o selectp2[75]
o selectp2[76]
o selectp2[77]
o selectp2[78]
o selectp2[79]
o selectp2[80]
o selectp2[81]
o selectp2[82]
o selectp2[83]
o selectp2[84]
o selectp2[85]
o selectp2[86]
o selectp2[87]
o selectp2[88]
o selectp2[89]
o selectp2[90]
o selectp2[91]
o selectp2[92]
o selectp2[93]
o selectp2[94]
o selectp2[95]
o selectp2[96]
o selectp2[97]
o selectp2[98]
o selectp2[99]
o selectp2[100]
o selectp2[101]
o selectp2[102]
o selectp2[103]
o selectp2[104]
o selectp2[105]
o selectp2[106]
o selectp2[107]
o selectp2[108]
o selectp2[109]
o selectp2[110]
o selectp2[111]
o selectp2[112]
o selectp2[113]
o selectp2[114]
o selectp2[115]
o selectp2[116]
o selectp2[117]
o selectp2[118]
o selectp2[119]
o selectp2[120]
o selectp2[121]
o selectp2[122]
o selectp2[123]
o selectp2[124]
o selectp2[125]
o selectp2[126]
o selectp2[127]
