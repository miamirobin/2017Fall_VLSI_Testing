name multi
i a[0]
i a[1]
i a[2]
i a[3]
i a[4]
i a[5]
i a[6]
i a[7]
i a[8]
i a[9]
i a[10]
i a[11]
i a[12]
i a[13]
i a[14]
i a[15]
i a[16]
i a[17]
i a[18]
i a[19]
i a[20]
i a[21]
i a[22]
i a[23]
i a[24]
i a[25]
i a[26]
i a[27]
i a[28]
i a[29]
i a[30]
i a[31]
i a[32]
i a[33]
i a[34]
i a[35]
i a[36]
i a[37]
i a[38]
i a[39]
i a[40]
i a[41]
i a[42]
i a[43]
i a[44]
i a[45]
i a[46]
i a[47]
i a[48]
i a[49]
i a[50]
i a[51]
i a[52]
i a[53]
i a[54]
i a[55]
i a[56]
i a[57]
i a[58]
i a[59]
i a[60]
i a[61]
i a[62]
i a[63]
i b[0]
i b[1]
i b[2]
i b[3]
i b[4]
i b[5]
i b[6]
i b[7]
i b[8]
i b[9]
i b[10]
i b[11]
i b[12]
i b[13]
i b[14]
i b[15]
i b[16]
i b[17]
i b[18]
i b[19]
i b[20]
i b[21]
i b[22]
i b[23]
i b[24]
i b[25]
i b[26]
i b[27]
i b[28]
i b[29]
i b[30]
i b[31]
i b[32]
i b[33]
i b[34]
i b[35]
i b[36]
i b[37]
i b[38]
i b[39]
i b[40]
i b[41]
i b[42]
i b[43]
i b[44]
i b[45]
i b[46]
i b[47]
i b[48]
i b[49]
i b[50]
i b[51]
i b[52]
i b[53]
i b[54]
i b[55]
i b[56]
i b[57]
i b[58]
i b[59]
i b[60]
i b[61]
i b[62]
i b[63]

g1 and a[0] b[0] ; n257
g2 and a[2] n257_not ; n258
g3 and a[2]_not n257_not ; n259
g4 and n258_not n259_not ; f[0]
g5 and a[0]_not a[1] ; n261
g6 and b[0] n261 ; n262
g7 and a[1]_not a[2] ; n263
g8 and a[1] a[2]_not ; n264
g9 and n263_not n264_not ; n265
g10 and a[0] n265 ; n266
g11 and b[1] n266 ; n267
g12 and n262_not n267_not ; n268
g13 and a[0] n265_not ; n269
g14 and b[0] b[1]_not ; n270
g15 and b[0]_not b[1] ; n271
g16 and n270_not n271_not ; n272
g17 and n269 n272_not ; n273
g18 and n268 n273_not ; n274
g19 and a[2] n274_not ; n275
g20 and a[2] n275_not ; n276
g21 and n274_not n275_not ; n277
g22 and n276_not n277_not ; n278
g23 and n258 n278_not ; n279
g24 and n258_not n278 ; n280
g25 and n279_not n280_not ; f[1]
g26 and b[2] n266 ; n282
g27 and a[0]_not n265_not ; n283
g28 and a[1]_not n283 ; n284
g29 and b[0] n284 ; n285
g30 and b[1] n261 ; n286
g31 and n285_not n286_not ; n287
g32 and n282_not n287 ; n288
g33 and b[0] b[2]_not ; n289
g34 and b[1] n289 ; n290
g35 and b[1] b[2]_not ; n291
g36 and b[1]_not b[2] ; n292
g37 and n291_not n292_not ; n293
g38 and b[0] b[1] ; n294
g39 and n293 n294_not ; n295
g40 and n290_not n295_not ; n296
g41 and n269 n296 ; n297
g42 and n288 n297_not ; n298
g43 and a[2] n298_not ; n299
g44 and a[2] n299_not ; n300
g45 and n298_not n299_not ; n301
g46 and n300_not n301_not ; n302
g47 and n279 n302_not ; n303
g48 and n279_not n302 ; n304
g49 and n303_not n304_not ; f[2]
g50 and b[3] n266 ; n306
g51 and b[1] n284 ; n307
g52 and b[2] n261 ; n308
g53 and n307_not n308_not ; n309
g54 and n306_not n309 ; n310
g55 and b[1] b[2] ; n311
g56 and n290_not n311_not ; n312
g57 and b[2]_not b[3]_not ; n313
g58 and b[2] b[3] ; n314
g59 and n313_not n314_not ; n315
g60 and n312_not n315 ; n316
g61 and n312 n315_not ; n317
g62 and n316_not n317_not ; n318
g63 and n269 n318 ; n319
g64 and n310 n319_not ; n320
g65 and a[2] n320_not ; n321
g66 and a[2] n321_not ; n322
g67 and n320_not n321_not ; n323
g68 and n322_not n323_not ; n324
g69 and a[2] a[3]_not ; n325
g70 and a[2]_not a[3] ; n326
g71 and n325_not n326_not ; n327
g72 and b[0] n327_not ; n328
g73 and n324_not n328 ; n329
g74 and n324 n328_not ; n330
g75 and n329_not n330_not ; n331
g76 and n303 n331 ; n332
g77 and n303_not n331_not ; n333
g78 and n332_not n333_not ; f[3]
g79 and b[4] n266 ; n335
g80 and b[2] n284 ; n336
g81 and b[3] n261 ; n337
g82 and n336_not n337_not ; n338
g83 and n335_not n338 ; n339
g84 and n314_not n316_not ; n340
g85 and b[3]_not b[4]_not ; n341
g86 and b[3] b[4] ; n342
g87 and n341_not n342_not ; n343
g88 and n340_not n343 ; n344
g89 and n340 n343_not ; n345
g90 and n344_not n345_not ; n346
g91 and n269 n346 ; n347
g92 and n339 n347_not ; n348
g93 and a[2] n348_not ; n349
g94 and a[2] n349_not ; n350
g95 and n348_not n349_not ; n351
g96 and n350_not n351_not ; n352
g97 and a[5] n328_not ; n353
g98 and a[3]_not a[4] ; n354
g99 and a[3] a[4]_not ; n355
g100 and n354_not n355_not ; n356
g101 and n327 n356_not ; n357
g102 and b[0] n357 ; n358
g103 and a[4]_not a[5] ; n359
g104 and a[4] a[5]_not ; n360
g105 and n359_not n360_not ; n361
g106 and n327_not n361 ; n362
g107 and b[1] n362 ; n363
g108 and n358_not n363_not ; n364
g109 and n327_not n361_not ; n365
g110 and n272_not n365 ; n366
g111 and n364 n366_not ; n367
g112 and a[5] n367_not ; n368
g113 and a[5] n368_not ; n369
g114 and n367_not n368_not ; n370
g115 and n369_not n370_not ; n371
g116 and n353 n371_not ; n372
g117 and n353_not n371 ; n373
g118 and n372_not n373_not ; n374
g119 and n352_not n374 ; n375
g120 and n374 n375_not ; n376
g121 and n352_not n375_not ; n377
g122 and n376_not n377_not ; n378
g123 and n329_not n332_not ; n379
g124 and n378_not n379_not ; n380
g125 and n378 n379 ; n381
g126 and n380_not n381_not ; f[4]
g127 and b[5] n266 ; n383
g128 and b[3] n284 ; n384
g129 and b[4] n261 ; n385
g130 and n384_not n385_not ; n386
g131 and n383_not n386 ; n387
g132 and n342_not n344_not ; n388
g133 and b[4]_not b[5]_not ; n389
g134 and b[4] b[5] ; n390
g135 and n389_not n390_not ; n391
g136 and n388_not n391 ; n392
g137 and n388 n391_not ; n393
g138 and n392_not n393_not ; n394
g139 and n269 n394 ; n395
g140 and n387 n395_not ; n396
g141 and a[2] n396_not ; n397
g142 and a[2] n397_not ; n398
g143 and n396_not n397_not ; n399
g144 and n398_not n399_not ; n400
g145 and b[2] n362 ; n401
g146 and n327 n361_not ; n402
g147 and n356 n402 ; n403
g148 and b[0] n403 ; n404
g149 and b[1] n357 ; n405
g150 and n404_not n405_not ; n406
g151 and n401_not n406 ; n407
g152 and n365_not n407 ; n408
g153 and n296_not n407 ; n409
g154 and n408_not n409_not ; n410
g155 and a[5] n410_not ; n411
g156 and a[5]_not n410 ; n412
g157 and n411_not n412_not ; n413
g158 and n372 n413_not ; n414
g159 and n372_not n413 ; n415
g160 and n414_not n415_not ; n416
g161 and n400_not n416 ; n417
g162 and n416 n417_not ; n418
g163 and n400_not n417_not ; n419
g164 and n418_not n419_not ; n420
g165 and n375_not n380_not ; n421
g166 and n420_not n421_not ; n422
g167 and n420 n421 ; n423
g168 and n422_not n423_not ; f[5]
g169 and n417_not n422_not ; n425
g170 and a[5] a[6]_not ; n426
g171 and a[5]_not a[6] ; n427
g172 and n426_not n427_not ; n428
g173 and b[0] n428_not ; n429
g174 and n414 n429 ; n430
g175 and n414 n430_not ; n431
g176 and n429 n430_not ; n432
g177 and n431_not n432_not ; n433
g178 and b[3] n362 ; n434
g179 and b[1] n403 ; n435
g180 and b[2] n357 ; n436
g181 and n435_not n436_not ; n437
g182 and n434_not n437 ; n438
g183 and n318 n365 ; n439
g184 and n438 n439_not ; n440
g185 and a[5] n440_not ; n441
g186 and a[5] n441_not ; n442
g187 and n440_not n441_not ; n443
g188 and n442_not n443_not ; n444
g189 and n433_not n444 ; n445
g190 and n433 n444_not ; n446
g191 and n445_not n446_not ; n447
g192 and b[6] n266 ; n448
g193 and b[4] n284 ; n449
g194 and b[5] n261 ; n450
g195 and n449_not n450_not ; n451
g196 and n448_not n451 ; n452
g197 and n390_not n392_not ; n453
g198 and b[5]_not b[6]_not ; n454
g199 and b[5] b[6] ; n455
g200 and n454_not n455_not ; n456
g201 and n453_not n456 ; n457
g202 and n453 n456_not ; n458
g203 and n457_not n458_not ; n459
g204 and n269 n459 ; n460
g205 and n452 n460_not ; n461
g206 and a[2] n461_not ; n462
g207 and a[2] n462_not ; n463
g208 and n461_not n462_not ; n464
g209 and n463_not n464_not ; n465
g210 and n447_not n465_not ; n466
g211 and n447 n465 ; n467
g212 and n466_not n467_not ; n468
g213 and n425_not n468 ; n469
g214 and n425 n468_not ; n470
g215 and n469_not n470_not ; f[6]
g216 and n466_not n469_not ; n472
g217 and b[7] n266 ; n473
g218 and b[5] n284 ; n474
g219 and b[6] n261 ; n475
g220 and n474_not n475_not ; n476
g221 and n473_not n476 ; n477
g222 and n455_not n457_not ; n478
g223 and b[6]_not b[7]_not ; n479
g224 and b[6] b[7] ; n480
g225 and n479_not n480_not ; n481
g226 and n478_not n481 ; n482
g227 and n478 n481_not ; n483
g228 and n482_not n483_not ; n484
g229 and n269 n484 ; n485
g230 and n477 n485_not ; n486
g231 and a[2] n486_not ; n487
g232 and a[2] n487_not ; n488
g233 and n486_not n487_not ; n489
g234 and n488_not n489_not ; n490
g235 and b[4] n362 ; n491
g236 and b[2] n403 ; n492
g237 and b[3] n357 ; n493
g238 and n492_not n493_not ; n494
g239 and n491_not n494 ; n495
g240 and n346 n365 ; n496
g241 and n495 n496_not ; n497
g242 and a[5] n497_not ; n498
g243 and a[5] n498_not ; n499
g244 and n497_not n498_not ; n500
g245 and n499_not n500_not ; n501
g246 and a[8] n429_not ; n502
g247 and a[6]_not a[7] ; n503
g248 and a[6] a[7]_not ; n504
g249 and n503_not n504_not ; n505
g250 and n428 n505_not ; n506
g251 and b[0] n506 ; n507
g252 and a[7]_not a[8] ; n508
g253 and a[7] a[8]_not ; n509
g254 and n508_not n509_not ; n510
g255 and n428_not n510 ; n511
g256 and b[1] n511 ; n512
g257 and n507_not n512_not ; n513
g258 and n428_not n510_not ; n514
g259 and n272_not n514 ; n515
g260 and n513 n515_not ; n516
g261 and a[8] n516_not ; n517
g262 and a[8] n517_not ; n518
g263 and n516_not n517_not ; n519
g264 and n518_not n519_not ; n520
g265 and n502 n520_not ; n521
g266 and n502_not n520 ; n522
g267 and n521_not n522_not ; n523
g268 and n501_not n523 ; n524
g269 and n523 n524_not ; n525
g270 and n501_not n524_not ; n526
g271 and n525_not n526_not ; n527
g272 and n433_not n444_not ; n528
g273 and n430_not n528_not ; n529
g274 and n527_not n529_not ; n530
g275 and n527 n529 ; n531
g276 and n530_not n531_not ; n532
g277 and n490_not n532 ; n533
g278 and n490 n532_not ; n534
g279 and n533_not n534_not ; n535
g280 and n472_not n535 ; n536
g281 and n472 n535_not ; n537
g282 and n536_not n537_not ; f[7]
g283 and b[2] n511 ; n539
g284 and n428 n510_not ; n540
g285 and n505 n540 ; n541
g286 and b[0] n541 ; n542
g287 and b[1] n506 ; n543
g288 and n542_not n543_not ; n544
g289 and n539_not n544 ; n545
g290 and n296 n514 ; n546
g291 and n545 n546_not ; n547
g292 and a[8] n547_not ; n548
g293 and a[8] n548_not ; n549
g294 and n547_not n548_not ; n550
g295 and n549_not n550_not ; n551
g296 and n521_not n551 ; n552
g297 and n521 n551_not ; n553
g298 and n552_not n553_not ; n554
g299 and b[5] n362 ; n555
g300 and b[3] n403 ; n556
g301 and b[4] n357 ; n557
g302 and n556_not n557_not ; n558
g303 and n555_not n558 ; n559
g304 and n365 n394 ; n560
g305 and n559 n560_not ; n561
g306 and a[5] n561_not ; n562
g307 and a[5] n562_not ; n563
g308 and n561_not n562_not ; n564
g309 and n563_not n564_not ; n565
g310 and n554 n565_not ; n566
g311 and n554 n566_not ; n567
g312 and n565_not n566_not ; n568
g313 and n567_not n568_not ; n569
g314 and n524_not n530_not ; n570
g315 and n569 n570 ; n571
g316 and n569_not n570_not ; n572
g317 and n571_not n572_not ; n573
g318 and b[8] n266 ; n574
g319 and b[6] n284 ; n575
g320 and b[7] n261 ; n576
g321 and n575_not n576_not ; n577
g322 and n574_not n577 ; n578
g323 and n480_not n482_not ; n579
g324 and b[7]_not b[8]_not ; n580
g325 and b[7] b[8] ; n581
g326 and n580_not n581_not ; n582
g327 and n579_not n582 ; n583
g328 and n579 n582_not ; n584
g329 and n583_not n584_not ; n585
g330 and n269 n585 ; n586
g331 and n578 n586_not ; n587
g332 and a[2] n587_not ; n588
g333 and a[2] n588_not ; n589
g334 and n587_not n588_not ; n590
g335 and n589_not n590_not ; n591
g336 and n573 n591_not ; n592
g337 and n573 n592_not ; n593
g338 and n591_not n592_not ; n594
g339 and n593_not n594_not ; n595
g340 and n533_not n536_not ; n596
g341 and n595_not n596_not ; n597
g342 and n595 n596 ; n598
g343 and n597_not n598_not ; f[8]
g344 and b[6] n362 ; n600
g345 and b[4] n403 ; n601
g346 and b[5] n357 ; n602
g347 and n601_not n602_not ; n603
g348 and n600_not n603 ; n604
g349 and n365 n459 ; n605
g350 and n604 n605_not ; n606
g351 and a[5] n606_not ; n607
g352 and a[5] n607_not ; n608
g353 and n606_not n607_not ; n609
g354 and n608_not n609_not ; n610
g355 and a[8] a[9]_not ; n611
g356 and a[8]_not a[9] ; n612
g357 and n611_not n612_not ; n613
g358 and b[0] n613_not ; n614
g359 and n553_not n614 ; n615
g360 and n553 n614_not ; n616
g361 and n615_not n616_not ; n617
g362 and b[3] n511 ; n618
g363 and b[1] n541 ; n619
g364 and b[2] n506 ; n620
g365 and n619_not n620_not ; n621
g366 and n618_not n621 ; n622
g367 and n318 n514 ; n623
g368 and n622 n623_not ; n624
g369 and a[8] n624_not ; n625
g370 and a[8] n625_not ; n626
g371 and n624_not n625_not ; n627
g372 and n626_not n627_not ; n628
g373 and n617_not n628_not ; n629
g374 and n617 n628 ; n630
g375 and n629_not n630_not ; n631
g376 and n610_not n631 ; n632
g377 and n631 n632_not ; n633
g378 and n610_not n632_not ; n634
g379 and n633_not n634_not ; n635
g380 and n566_not n572_not ; n636
g381 and n635 n636 ; n637
g382 and n635_not n636_not ; n638
g383 and n637_not n638_not ; n639
g384 and b[9] n266 ; n640
g385 and b[7] n284 ; n641
g386 and b[8] n261 ; n642
g387 and n641_not n642_not ; n643
g388 and n640_not n643 ; n644
g389 and n581_not n583_not ; n645
g390 and b[8]_not b[9]_not ; n646
g391 and b[8] b[9] ; n647
g392 and n646_not n647_not ; n648
g393 and n645_not n648 ; n649
g394 and n645 n648_not ; n650
g395 and n649_not n650_not ; n651
g396 and n269 n651 ; n652
g397 and n644 n652_not ; n653
g398 and a[2] n653_not ; n654
g399 and a[2] n654_not ; n655
g400 and n653_not n654_not ; n656
g401 and n655_not n656_not ; n657
g402 and n639 n657_not ; n658
g403 and n639 n658_not ; n659
g404 and n657_not n658_not ; n660
g405 and n659_not n660_not ; n661
g406 and n592_not n597_not ; n662
g407 and n661_not n662_not ; n663
g408 and n661 n662 ; n664
g409 and n663_not n664_not ; f[9]
g410 and n658_not n663_not ; n666
g411 and b[7] n362 ; n667
g412 and b[5] n403 ; n668
g413 and b[6] n357 ; n669
g414 and n668_not n669_not ; n670
g415 and n667_not n670 ; n671
g416 and n365 n484 ; n672
g417 and n671 n672_not ; n673
g418 and a[5] n673_not ; n674
g419 and a[5] n674_not ; n675
g420 and n673_not n674_not ; n676
g421 and n675_not n676_not ; n677
g422 and n553 n614 ; n678
g423 and n629_not n678_not ; n679
g424 and b[4] n511 ; n680
g425 and b[2] n541 ; n681
g426 and b[3] n506 ; n682
g427 and n681_not n682_not ; n683
g428 and n680_not n683 ; n684
g429 and n346 n514 ; n685
g430 and n684 n685_not ; n686
g431 and a[8] n686_not ; n687
g432 and a[8] n687_not ; n688
g433 and n686_not n687_not ; n689
g434 and n688_not n689_not ; n690
g435 and a[11] n614_not ; n691
g436 and a[9]_not a[10] ; n692
g437 and a[9] a[10]_not ; n693
g438 and n692_not n693_not ; n694
g439 and n613 n694_not ; n695
g440 and b[0] n695 ; n696
g441 and a[10]_not a[11] ; n697
g442 and a[10] a[11]_not ; n698
g443 and n697_not n698_not ; n699
g444 and n613_not n699 ; n700
g445 and b[1] n700 ; n701
g446 and n696_not n701_not ; n702
g447 and n613_not n699_not ; n703
g448 and n272_not n703 ; n704
g449 and n702 n704_not ; n705
g450 and a[11] n705_not ; n706
g451 and a[11] n706_not ; n707
g452 and n705_not n706_not ; n708
g453 and n707_not n708_not ; n709
g454 and n691 n709_not ; n710
g455 and n691_not n709 ; n711
g456 and n710_not n711_not ; n712
g457 and n690 n712_not ; n713
g458 and n690_not n712 ; n714
g459 and n713_not n714_not ; n715
g460 and n679_not n715 ; n716
g461 and n679 n715_not ; n717
g462 and n716_not n717_not ; n718
g463 and n677_not n718 ; n719
g464 and n718 n719_not ; n720
g465 and n677_not n719_not ; n721
g466 and n720_not n721_not ; n722
g467 and n632_not n638_not ; n723
g468 and n722 n723 ; n724
g469 and n722_not n723_not ; n725
g470 and n724_not n725_not ; n726
g471 and b[10] n266 ; n727
g472 and b[8] n284 ; n728
g473 and b[9] n261 ; n729
g474 and n728_not n729_not ; n730
g475 and n727_not n730 ; n731
g476 and n647_not n649_not ; n732
g477 and b[9]_not b[10]_not ; n733
g478 and b[9] b[10] ; n734
g479 and n733_not n734_not ; n735
g480 and n732_not n735 ; n736
g481 and n732 n735_not ; n737
g482 and n736_not n737_not ; n738
g483 and n269 n738 ; n739
g484 and n731 n739_not ; n740
g485 and a[2] n740_not ; n741
g486 and a[2] n741_not ; n742
g487 and n740_not n741_not ; n743
g488 and n742_not n743_not ; n744
g489 and n726_not n744 ; n745
g490 and n726 n744_not ; n746
g491 and n745_not n746_not ; n747
g492 and n666_not n747 ; n748
g493 and n666 n747_not ; n749
g494 and n748_not n749_not ; f[10]
g495 and n746_not n748_not ; n751
g496 and n719_not n725_not ; n752
g497 and b[8] n362 ; n753
g498 and b[6] n403 ; n754
g499 and b[7] n357 ; n755
g500 and n754_not n755_not ; n756
g501 and n753_not n756 ; n757
g502 and n365 n585 ; n758
g503 and n757 n758_not ; n759
g504 and a[5] n759_not ; n760
g505 and a[5] n760_not ; n761
g506 and n759_not n760_not ; n762
g507 and n761_not n762_not ; n763
g508 and n714_not n716_not ; n764
g509 and b[2] n700 ; n765
g510 and n613 n699_not ; n766
g511 and n694 n766 ; n767
g512 and b[0] n767 ; n768
g513 and b[1] n695 ; n769
g514 and n768_not n769_not ; n770
g515 and n765_not n770 ; n771
g516 and n296 n703 ; n772
g517 and n771 n772_not ; n773
g518 and a[11] n773_not ; n774
g519 and a[11] n774_not ; n775
g520 and n773_not n774_not ; n776
g521 and n775_not n776_not ; n777
g522 and n710_not n777 ; n778
g523 and n710 n777_not ; n779
g524 and n778_not n779_not ; n780
g525 and b[5] n511 ; n781
g526 and b[3] n541 ; n782
g527 and b[4] n506 ; n783
g528 and n782_not n783_not ; n784
g529 and n781_not n784 ; n785
g530 and n394 n514 ; n786
g531 and n785 n786_not ; n787
g532 and a[8] n787_not ; n788
g533 and a[8] n788_not ; n789
g534 and n787_not n788_not ; n790
g535 and n789_not n790_not ; n791
g536 and n780 n791_not ; n792
g537 and n780 n792_not ; n793
g538 and n791_not n792_not ; n794
g539 and n793_not n794_not ; n795
g540 and n764_not n795_not ; n796
g541 and n764 n795 ; n797
g542 and n796_not n797_not ; n798
g543 and n763_not n798 ; n799
g544 and n763_not n799_not ; n800
g545 and n798 n799_not ; n801
g546 and n800_not n801_not ; n802
g547 and n752_not n802_not ; n803
g548 and n752_not n803_not ; n804
g549 and n802_not n803_not ; n805
g550 and n804_not n805_not ; n806
g551 and b[11] n266 ; n807
g552 and b[9] n284 ; n808
g553 and b[10] n261 ; n809
g554 and n808_not n809_not ; n810
g555 and n807_not n810 ; n811
g556 and n734_not n736_not ; n812
g557 and b[10]_not b[11]_not ; n813
g558 and b[10] b[11] ; n814
g559 and n813_not n814_not ; n815
g560 and n812_not n815 ; n816
g561 and n812 n815_not ; n817
g562 and n816_not n817_not ; n818
g563 and n269 n818 ; n819
g564 and n811 n819_not ; n820
g565 and a[2] n820_not ; n821
g566 and a[2] n821_not ; n822
g567 and n820_not n821_not ; n823
g568 and n822_not n823_not ; n824
g569 and n806_not n824 ; n825
g570 and n806 n824_not ; n826
g571 and n825_not n826_not ; n827
g572 and n751_not n827_not ; n828
g573 and n751 n827 ; n829
g574 and n828_not n829_not ; f[11]
g575 and b[12] n266 ; n831
g576 and b[10] n284 ; n832
g577 and b[11] n261 ; n833
g578 and n832_not n833_not ; n834
g579 and n831_not n834 ; n835
g580 and n814_not n816_not ; n836
g581 and b[11]_not b[12]_not ; n837
g582 and b[11] b[12] ; n838
g583 and n837_not n838_not ; n839
g584 and n836_not n839 ; n840
g585 and n836 n839_not ; n841
g586 and n840_not n841_not ; n842
g587 and n269 n842 ; n843
g588 and n835 n843_not ; n844
g589 and a[2] n844_not ; n845
g590 and a[2] n845_not ; n846
g591 and n844_not n845_not ; n847
g592 and n846_not n847_not ; n848
g593 and b[6] n511 ; n849
g594 and b[4] n541 ; n850
g595 and b[5] n506 ; n851
g596 and n850_not n851_not ; n852
g597 and n849_not n852 ; n853
g598 and n459 n514 ; n854
g599 and n853 n854_not ; n855
g600 and a[8] n855_not ; n856
g601 and a[8] n856_not ; n857
g602 and n855_not n856_not ; n858
g603 and n857_not n858_not ; n859
g604 and a[11] a[12]_not ; n860
g605 and a[11]_not a[12] ; n861
g606 and n860_not n861_not ; n862
g607 and b[0] n862_not ; n863
g608 and n779_not n863 ; n864
g609 and n779 n863_not ; n865
g610 and n864_not n865_not ; n866
g611 and b[3] n700 ; n867
g612 and b[1] n767 ; n868
g613 and b[2] n695 ; n869
g614 and n868_not n869_not ; n870
g615 and n867_not n870 ; n871
g616 and n318 n703 ; n872
g617 and n871 n872_not ; n873
g618 and a[11] n873_not ; n874
g619 and a[11] n874_not ; n875
g620 and n873_not n874_not ; n876
g621 and n875_not n876_not ; n877
g622 and n866_not n877_not ; n878
g623 and n866 n877 ; n879
g624 and n878_not n879_not ; n880
g625 and n859_not n880 ; n881
g626 and n880 n881_not ; n882
g627 and n859_not n881_not ; n883
g628 and n882_not n883_not ; n884
g629 and n792_not n796_not ; n885
g630 and n884 n885 ; n886
g631 and n884_not n885_not ; n887
g632 and n886_not n887_not ; n888
g633 and b[9] n362 ; n889
g634 and b[7] n403 ; n890
g635 and b[8] n357 ; n891
g636 and n890_not n891_not ; n892
g637 and n889_not n892 ; n893
g638 and n365 n651 ; n894
g639 and n893 n894_not ; n895
g640 and a[5] n895_not ; n896
g641 and a[5] n896_not ; n897
g642 and n895_not n896_not ; n898
g643 and n897_not n898_not ; n899
g644 and n888_not n899 ; n900
g645 and n888 n899_not ; n901
g646 and n900_not n901_not ; n902
g647 and n799_not n803_not ; n903
g648 and n902 n903_not ; n904
g649 and n902_not n903 ; n905
g650 and n904_not n905_not ; n906
g651 and n848_not n906 ; n907
g652 and n906 n907_not ; n908
g653 and n848_not n907_not ; n909
g654 and n908_not n909_not ; n910
g655 and n806_not n824_not ; n911
g656 and n828_not n911_not ; n912
g657 and n910_not n912_not ; n913
g658 and n910 n912 ; n914
g659 and n913_not n914_not ; f[12]
g660 and n907_not n913_not ; n916
g661 and n901_not n904_not ; n917
g662 and b[7] n511 ; n918
g663 and b[5] n541 ; n919
g664 and b[6] n506 ; n920
g665 and n919_not n920_not ; n921
g666 and n918_not n921 ; n922
g667 and n484 n514 ; n923
g668 and n922 n923_not ; n924
g669 and a[8] n924_not ; n925
g670 and a[8] n925_not ; n926
g671 and n924_not n925_not ; n927
g672 and n926_not n927_not ; n928
g673 and n779 n863 ; n929
g674 and n878_not n929_not ; n930
g675 and b[4] n700 ; n931
g676 and b[2] n767 ; n932
g677 and b[3] n695 ; n933
g678 and n932_not n933_not ; n934
g679 and n931_not n934 ; n935
g680 and n346 n703 ; n936
g681 and n935 n936_not ; n937
g682 and a[11] n937_not ; n938
g683 and a[11] n938_not ; n939
g684 and n937_not n938_not ; n940
g685 and n939_not n940_not ; n941
g686 and a[14] n863_not ; n942
g687 and a[12]_not a[13] ; n943
g688 and a[12] a[13]_not ; n944
g689 and n943_not n944_not ; n945
g690 and n862 n945_not ; n946
g691 and b[0] n946 ; n947
g692 and a[13]_not a[14] ; n948
g693 and a[13] a[14]_not ; n949
g694 and n948_not n949_not ; n950
g695 and n862_not n950 ; n951
g696 and b[1] n951 ; n952
g697 and n947_not n952_not ; n953
g698 and n862_not n950_not ; n954
g699 and n272_not n954 ; n955
g700 and n953 n955_not ; n956
g701 and a[14] n956_not ; n957
g702 and a[14] n957_not ; n958
g703 and n956_not n957_not ; n959
g704 and n958_not n959_not ; n960
g705 and n942 n960_not ; n961
g706 and n942_not n960 ; n962
g707 and n961_not n962_not ; n963
g708 and n941 n963_not ; n964
g709 and n941_not n963 ; n965
g710 and n964_not n965_not ; n966
g711 and n930_not n966 ; n967
g712 and n930 n966_not ; n968
g713 and n967_not n968_not ; n969
g714 and n928_not n969 ; n970
g715 and n969 n970_not ; n971
g716 and n928_not n970_not ; n972
g717 and n971_not n972_not ; n973
g718 and n881_not n887_not ; n974
g719 and n973 n974 ; n975
g720 and n973_not n974_not ; n976
g721 and n975_not n976_not ; n977
g722 and b[10] n362 ; n978
g723 and b[8] n403 ; n979
g724 and b[9] n357 ; n980
g725 and n979_not n980_not ; n981
g726 and n978_not n981 ; n982
g727 and n365 n738 ; n983
g728 and n982 n983_not ; n984
g729 and a[5] n984_not ; n985
g730 and a[5] n985_not ; n986
g731 and n984_not n985_not ; n987
g732 and n986_not n987_not ; n988
g733 and n977 n988_not ; n989
g734 and n977_not n988 ; n990
g735 and n917_not n990_not ; n991
g736 and n989_not n991 ; n992
g737 and n917_not n992_not ; n993
g738 and n989_not n992_not ; n994
g739 and n990_not n994 ; n995
g740 and n993_not n995_not ; n996
g741 and b[13] n266 ; n997
g742 and b[11] n284 ; n998
g743 and b[12] n261 ; n999
g744 and n998_not n999_not ; n1000
g745 and n997_not n1000 ; n1001
g746 and n838_not n840_not ; n1002
g747 and b[12]_not b[13]_not ; n1003
g748 and b[12] b[13] ; n1004
g749 and n1003_not n1004_not ; n1005
g750 and n1002_not n1005 ; n1006
g751 and n1002 n1005_not ; n1007
g752 and n1006_not n1007_not ; n1008
g753 and n269 n1008 ; n1009
g754 and n1001 n1009_not ; n1010
g755 and a[2] n1010_not ; n1011
g756 and a[2] n1011_not ; n1012
g757 and n1010_not n1011_not ; n1013
g758 and n1012_not n1013_not ; n1014
g759 and n996_not n1014 ; n1015
g760 and n996 n1014_not ; n1016
g761 and n1015_not n1016_not ; n1017
g762 and n916_not n1017_not ; n1018
g763 and n916 n1017 ; n1019
g764 and n1018_not n1019_not ; f[13]
g765 and n996_not n1014_not ; n1021
g766 and n1018_not n1021_not ; n1022
g767 and b[14] n266 ; n1023
g768 and b[12] n284 ; n1024
g769 and b[13] n261 ; n1025
g770 and n1024_not n1025_not ; n1026
g771 and n1023_not n1026 ; n1027
g772 and n1004_not n1006_not ; n1028
g773 and b[13]_not b[14]_not ; n1029
g774 and b[13] b[14] ; n1030
g775 and n1029_not n1030_not ; n1031
g776 and n1028_not n1031 ; n1032
g777 and n1028 n1031_not ; n1033
g778 and n1032_not n1033_not ; n1034
g779 and n269 n1034 ; n1035
g780 and n1027 n1035_not ; n1036
g781 and a[2] n1036_not ; n1037
g782 and a[2] n1037_not ; n1038
g783 and n1036_not n1037_not ; n1039
g784 and n1038_not n1039_not ; n1040
g785 and b[11] n362 ; n1041
g786 and b[9] n403 ; n1042
g787 and b[10] n357 ; n1043
g788 and n1042_not n1043_not ; n1044
g789 and n1041_not n1044 ; n1045
g790 and n365 n818 ; n1046
g791 and n1045 n1046_not ; n1047
g792 and a[5] n1047_not ; n1048
g793 and a[5] n1048_not ; n1049
g794 and n1047_not n1048_not ; n1050
g795 and n1049_not n1050_not ; n1051
g796 and n970_not n976_not ; n1052
g797 and n965_not n967_not ; n1053
g798 and b[2] n951 ; n1054
g799 and n862 n950_not ; n1055
g800 and n945 n1055 ; n1056
g801 and b[0] n1056 ; n1057
g802 and b[1] n946 ; n1058
g803 and n1057_not n1058_not ; n1059
g804 and n1054_not n1059 ; n1060
g805 and n296 n954 ; n1061
g806 and n1060 n1061_not ; n1062
g807 and a[14] n1062_not ; n1063
g808 and a[14] n1063_not ; n1064
g809 and n1062_not n1063_not ; n1065
g810 and n1064_not n1065_not ; n1066
g811 and n961_not n1066 ; n1067
g812 and n961 n1066_not ; n1068
g813 and n1067_not n1068_not ; n1069
g814 and b[5] n700 ; n1070
g815 and b[3] n767 ; n1071
g816 and b[4] n695 ; n1072
g817 and n1071_not n1072_not ; n1073
g818 and n1070_not n1073 ; n1074
g819 and n394 n703 ; n1075
g820 and n1074 n1075_not ; n1076
g821 and a[11] n1076_not ; n1077
g822 and a[11] n1077_not ; n1078
g823 and n1076_not n1077_not ; n1079
g824 and n1078_not n1079_not ; n1080
g825 and n1069 n1080_not ; n1081
g826 and n1069_not n1080 ; n1082
g827 and n1053_not n1082_not ; n1083
g828 and n1081_not n1083 ; n1084
g829 and n1053_not n1084_not ; n1085
g830 and n1081_not n1084_not ; n1086
g831 and n1082_not n1086 ; n1087
g832 and n1085_not n1087_not ; n1088
g833 and b[8] n511 ; n1089
g834 and b[6] n541 ; n1090
g835 and b[7] n506 ; n1091
g836 and n1090_not n1091_not ; n1092
g837 and n1089_not n1092 ; n1093
g838 and n514 n585 ; n1094
g839 and n1093 n1094_not ; n1095
g840 and a[8] n1095_not ; n1096
g841 and a[8] n1096_not ; n1097
g842 and n1095_not n1096_not ; n1098
g843 and n1097_not n1098_not ; n1099
g844 and n1088 n1099 ; n1100
g845 and n1088_not n1099_not ; n1101
g846 and n1100_not n1101_not ; n1102
g847 and n1052_not n1102 ; n1103
g848 and n1052 n1102_not ; n1104
g849 and n1103_not n1104_not ; n1105
g850 and n1051 n1105_not ; n1106
g851 and n1051_not n1105 ; n1107
g852 and n1106_not n1107_not ; n1108
g853 and n994_not n1108 ; n1109
g854 and n994 n1108_not ; n1110
g855 and n1109_not n1110_not ; n1111
g856 and n1040 n1111 ; n1112
g857 and n1040_not n1111_not ; n1113
g858 and n1112_not n1113_not ; n1114
g859 and n1022_not n1114_not ; n1115
g860 and n1022 n1114 ; n1116
g861 and n1115_not n1116_not ; f[14]
g862 and n1040_not n1111 ; n1118
g863 and n1115_not n1118_not ; n1119
g864 and b[15] n266 ; n1120
g865 and b[13] n284 ; n1121
g866 and b[14] n261 ; n1122
g867 and n1121_not n1122_not ; n1123
g868 and n1120_not n1123 ; n1124
g869 and n1030_not n1032_not ; n1125
g870 and b[14]_not b[15]_not ; n1126
g871 and b[14] b[15] ; n1127
g872 and n1126_not n1127_not ; n1128
g873 and n1125_not n1128 ; n1129
g874 and n1125 n1128_not ; n1130
g875 and n1129_not n1130_not ; n1131
g876 and n269 n1131 ; n1132
g877 and n1124 n1132_not ; n1133
g878 and a[2] n1133_not ; n1134
g879 and a[2] n1134_not ; n1135
g880 and n1133_not n1134_not ; n1136
g881 and n1135_not n1136_not ; n1137
g882 and n1107_not n1109_not ; n1138
g883 and b[12] n362 ; n1139
g884 and b[10] n403 ; n1140
g885 and b[11] n357 ; n1141
g886 and n1140_not n1141_not ; n1142
g887 and n1139_not n1142 ; n1143
g888 and n365 n842 ; n1144
g889 and n1143 n1144_not ; n1145
g890 and a[5] n1145_not ; n1146
g891 and a[5] n1146_not ; n1147
g892 and n1145_not n1146_not ; n1148
g893 and n1147_not n1148_not ; n1149
g894 and n1101_not n1103_not ; n1150
g895 and b[9] n511 ; n1151
g896 and b[7] n541 ; n1152
g897 and b[8] n506 ; n1153
g898 and n1152_not n1153_not ; n1154
g899 and n1151_not n1154 ; n1155
g900 and n514 n651 ; n1156
g901 and n1155 n1156_not ; n1157
g902 and a[8] n1157_not ; n1158
g903 and a[8] n1158_not ; n1159
g904 and n1157_not n1158_not ; n1160
g905 and n1159_not n1160_not ; n1161
g906 and b[6] n700 ; n1162
g907 and b[4] n767 ; n1163
g908 and b[5] n695 ; n1164
g909 and n1163_not n1164_not ; n1165
g910 and n1162_not n1165 ; n1166
g911 and n459 n703 ; n1167
g912 and n1166 n1167_not ; n1168
g913 and a[11] n1168_not ; n1169
g914 and a[11] n1169_not ; n1170
g915 and n1168_not n1169_not ; n1171
g916 and n1170_not n1171_not ; n1172
g917 and a[14] a[15]_not ; n1173
g918 and a[14]_not a[15] ; n1174
g919 and n1173_not n1174_not ; n1175
g920 and b[0] n1175_not ; n1176
g921 and n1068_not n1176 ; n1177
g922 and n1068 n1176_not ; n1178
g923 and n1177_not n1178_not ; n1179
g924 and b[3] n951 ; n1180
g925 and b[1] n1056 ; n1181
g926 and b[2] n946 ; n1182
g927 and n1181_not n1182_not ; n1183
g928 and n1180_not n1183 ; n1184
g929 and n318 n954 ; n1185
g930 and n1184 n1185_not ; n1186
g931 and a[14] n1186_not ; n1187
g932 and a[14] n1187_not ; n1188
g933 and n1186_not n1187_not ; n1189
g934 and n1188_not n1189_not ; n1190
g935 and n1179_not n1190_not ; n1191
g936 and n1179 n1190 ; n1192
g937 and n1191_not n1192_not ; n1193
g938 and n1172_not n1193 ; n1194
g939 and n1193 n1194_not ; n1195
g940 and n1172_not n1194_not ; n1196
g941 and n1195_not n1196_not ; n1197
g942 and n1086_not n1197_not ; n1198
g943 and n1086 n1197 ; n1199
g944 and n1198_not n1199_not ; n1200
g945 and n1161_not n1200 ; n1201
g946 and n1161_not n1201_not ; n1202
g947 and n1200 n1201_not ; n1203
g948 and n1202_not n1203_not ; n1204
g949 and n1150_not n1204_not ; n1205
g950 and n1150 n1203_not ; n1206
g951 and n1202_not n1206 ; n1207
g952 and n1205_not n1207_not ; n1208
g953 and n1149_not n1208 ; n1209
g954 and n1149_not n1209_not ; n1210
g955 and n1208 n1209_not ; n1211
g956 and n1210_not n1211_not ; n1212
g957 and n1138_not n1212_not ; n1213
g958 and n1138 n1211_not ; n1214
g959 and n1210_not n1214 ; n1215
g960 and n1213_not n1215_not ; n1216
g961 and n1137_not n1216 ; n1217
g962 and n1137_not n1217_not ; n1218
g963 and n1216 n1217_not ; n1219
g964 and n1218_not n1219_not ; n1220
g965 and n1119_not n1220_not ; n1221
g966 and n1119 n1219_not ; n1222
g967 and n1218_not n1222 ; n1223
g968 and n1221_not n1223_not ; f[15]
g969 and n1217_not n1221_not ; n1225
g970 and b[16] n266 ; n1226
g971 and b[14] n284 ; n1227
g972 and b[15] n261 ; n1228
g973 and n1227_not n1228_not ; n1229
g974 and n1226_not n1229 ; n1230
g975 and n1127_not n1129_not ; n1231
g976 and b[15]_not b[16]_not ; n1232
g977 and b[15] b[16] ; n1233
g978 and n1232_not n1233_not ; n1234
g979 and n1231_not n1234 ; n1235
g980 and n1231 n1234_not ; n1236
g981 and n1235_not n1236_not ; n1237
g982 and n269 n1237 ; n1238
g983 and n1230 n1238_not ; n1239
g984 and a[2] n1239_not ; n1240
g985 and a[2] n1240_not ; n1241
g986 and n1239_not n1240_not ; n1242
g987 and n1241_not n1242_not ; n1243
g988 and n1209_not n1213_not ; n1244
g989 and b[13] n362 ; n1245
g990 and b[11] n403 ; n1246
g991 and b[12] n357 ; n1247
g992 and n1246_not n1247_not ; n1248
g993 and n1245_not n1248 ; n1249
g994 and n365 n1008 ; n1250
g995 and n1249 n1250_not ; n1251
g996 and a[5] n1251_not ; n1252
g997 and a[5] n1252_not ; n1253
g998 and n1251_not n1252_not ; n1254
g999 and n1253_not n1254_not ; n1255
g1000 and n1201_not n1205_not ; n1256
g1001 and b[10] n511 ; n1257
g1002 and b[8] n541 ; n1258
g1003 and b[9] n506 ; n1259
g1004 and n1258_not n1259_not ; n1260
g1005 and n1257_not n1260 ; n1261
g1006 and n514 n738 ; n1262
g1007 and n1261 n1262_not ; n1263
g1008 and a[8] n1263_not ; n1264
g1009 and a[8] n1264_not ; n1265
g1010 and n1263_not n1264_not ; n1266
g1011 and n1265_not n1266_not ; n1267
g1012 and n1194_not n1198_not ; n1268
g1013 and b[7] n700 ; n1269
g1014 and b[5] n767 ; n1270
g1015 and b[6] n695 ; n1271
g1016 and n1270_not n1271_not ; n1272
g1017 and n1269_not n1272 ; n1273
g1018 and n484 n703 ; n1274
g1019 and n1273 n1274_not ; n1275
g1020 and a[11] n1275_not ; n1276
g1021 and a[11] n1276_not ; n1277
g1022 and n1275_not n1276_not ; n1278
g1023 and n1277_not n1278_not ; n1279
g1024 and n1068 n1176 ; n1280
g1025 and n1191_not n1280_not ; n1281
g1026 and b[4] n951 ; n1282
g1027 and b[2] n1056 ; n1283
g1028 and b[3] n946 ; n1284
g1029 and n1283_not n1284_not ; n1285
g1030 and n1282_not n1285 ; n1286
g1031 and n346 n954 ; n1287
g1032 and n1286 n1287_not ; n1288
g1033 and a[14] n1288_not ; n1289
g1034 and a[14] n1289_not ; n1290
g1035 and n1288_not n1289_not ; n1291
g1036 and n1290_not n1291_not ; n1292
g1037 and a[17] n1176_not ; n1293
g1038 and a[15]_not a[16] ; n1294
g1039 and a[15] a[16]_not ; n1295
g1040 and n1294_not n1295_not ; n1296
g1041 and n1175 n1296_not ; n1297
g1042 and b[0] n1297 ; n1298
g1043 and a[16]_not a[17] ; n1299
g1044 and a[16] a[17]_not ; n1300
g1045 and n1299_not n1300_not ; n1301
g1046 and n1175_not n1301 ; n1302
g1047 and b[1] n1302 ; n1303
g1048 and n1298_not n1303_not ; n1304
g1049 and n1175_not n1301_not ; n1305
g1050 and n272_not n1305 ; n1306
g1051 and n1304 n1306_not ; n1307
g1052 and a[17] n1307_not ; n1308
g1053 and a[17] n1308_not ; n1309
g1054 and n1307_not n1308_not ; n1310
g1055 and n1309_not n1310_not ; n1311
g1056 and n1293 n1311_not ; n1312
g1057 and n1293_not n1311 ; n1313
g1058 and n1312_not n1313_not ; n1314
g1059 and n1292 n1314_not ; n1315
g1060 and n1292_not n1314 ; n1316
g1061 and n1315_not n1316_not ; n1317
g1062 and n1281_not n1317 ; n1318
g1063 and n1281 n1317_not ; n1319
g1064 and n1318_not n1319_not ; n1320
g1065 and n1279 n1320_not ; n1321
g1066 and n1279_not n1320 ; n1322
g1067 and n1321_not n1322_not ; n1323
g1068 and n1268_not n1323 ; n1324
g1069 and n1268 n1323_not ; n1325
g1070 and n1324_not n1325_not ; n1326
g1071 and n1267 n1326_not ; n1327
g1072 and n1267_not n1326 ; n1328
g1073 and n1327_not n1328_not ; n1329
g1074 and n1256_not n1329 ; n1330
g1075 and n1256 n1329_not ; n1331
g1076 and n1330_not n1331_not ; n1332
g1077 and n1255 n1332_not ; n1333
g1078 and n1255_not n1332 ; n1334
g1079 and n1333_not n1334_not ; n1335
g1080 and n1244_not n1335 ; n1336
g1081 and n1244 n1335_not ; n1337
g1082 and n1336_not n1337_not ; n1338
g1083 and n1243 n1338 ; n1339
g1084 and n1243_not n1338_not ; n1340
g1085 and n1339_not n1340_not ; n1341
g1086 and n1225_not n1341_not ; n1342
g1087 and n1225 n1341 ; n1343
g1088 and n1342_not n1343_not ; f[16]
g1089 and b[17] n266 ; n1345
g1090 and b[15] n284 ; n1346
g1091 and b[16] n261 ; n1347
g1092 and n1346_not n1347_not ; n1348
g1093 and n1345_not n1348 ; n1349
g1094 and n1233_not n1235_not ; n1350
g1095 and b[16]_not b[17]_not ; n1351
g1096 and b[16] b[17] ; n1352
g1097 and n1351_not n1352_not ; n1353
g1098 and n1350_not n1353 ; n1354
g1099 and n1350 n1353_not ; n1355
g1100 and n1354_not n1355_not ; n1356
g1101 and n269 n1356 ; n1357
g1102 and n1349 n1357_not ; n1358
g1103 and a[2] n1358_not ; n1359
g1104 and a[2] n1359_not ; n1360
g1105 and n1358_not n1359_not ; n1361
g1106 and n1360_not n1361_not ; n1362
g1107 and n1334_not n1336_not ; n1363
g1108 and b[14] n362 ; n1364
g1109 and b[12] n403 ; n1365
g1110 and b[13] n357 ; n1366
g1111 and n1365_not n1366_not ; n1367
g1112 and n1364_not n1367 ; n1368
g1113 and n365 n1034 ; n1369
g1114 and n1368 n1369_not ; n1370
g1115 and a[5] n1370_not ; n1371
g1116 and a[5] n1371_not ; n1372
g1117 and n1370_not n1371_not ; n1373
g1118 and n1372_not n1373_not ; n1374
g1119 and n1328_not n1330_not ; n1375
g1120 and b[11] n511 ; n1376
g1121 and b[9] n541 ; n1377
g1122 and b[10] n506 ; n1378
g1123 and n1377_not n1378_not ; n1379
g1124 and n1376_not n1379 ; n1380
g1125 and n514 n818 ; n1381
g1126 and n1380 n1381_not ; n1382
g1127 and a[8] n1382_not ; n1383
g1128 and a[8] n1383_not ; n1384
g1129 and n1382_not n1383_not ; n1385
g1130 and n1384_not n1385_not ; n1386
g1131 and n1322_not n1324_not ; n1387
g1132 and n1316_not n1318_not ; n1388
g1133 and b[2] n1302 ; n1389
g1134 and n1175 n1301_not ; n1390
g1135 and n1296 n1390 ; n1391
g1136 and b[0] n1391 ; n1392
g1137 and b[1] n1297 ; n1393
g1138 and n1392_not n1393_not ; n1394
g1139 and n1389_not n1394 ; n1395
g1140 and n296 n1305 ; n1396
g1141 and n1395 n1396_not ; n1397
g1142 and a[17] n1397_not ; n1398
g1143 and a[17] n1398_not ; n1399
g1144 and n1397_not n1398_not ; n1400
g1145 and n1399_not n1400_not ; n1401
g1146 and n1312_not n1401 ; n1402
g1147 and n1312 n1401_not ; n1403
g1148 and n1402_not n1403_not ; n1404
g1149 and b[5] n951 ; n1405
g1150 and b[3] n1056 ; n1406
g1151 and b[4] n946 ; n1407
g1152 and n1406_not n1407_not ; n1408
g1153 and n1405_not n1408 ; n1409
g1154 and n394 n954 ; n1410
g1155 and n1409 n1410_not ; n1411
g1156 and a[14] n1411_not ; n1412
g1157 and a[14] n1412_not ; n1413
g1158 and n1411_not n1412_not ; n1414
g1159 and n1413_not n1414_not ; n1415
g1160 and n1404 n1415_not ; n1416
g1161 and n1404_not n1415 ; n1417
g1162 and n1388_not n1417_not ; n1418
g1163 and n1416_not n1418 ; n1419
g1164 and n1388_not n1419_not ; n1420
g1165 and n1416_not n1419_not ; n1421
g1166 and n1417_not n1421 ; n1422
g1167 and n1420_not n1422_not ; n1423
g1168 and b[8] n700 ; n1424
g1169 and b[6] n767 ; n1425
g1170 and b[7] n695 ; n1426
g1171 and n1425_not n1426_not ; n1427
g1172 and n1424_not n1427 ; n1428
g1173 and n585 n703 ; n1429
g1174 and n1428 n1429_not ; n1430
g1175 and a[11] n1430_not ; n1431
g1176 and a[11] n1431_not ; n1432
g1177 and n1430_not n1431_not ; n1433
g1178 and n1432_not n1433_not ; n1434
g1179 and n1423 n1434 ; n1435
g1180 and n1423_not n1434_not ; n1436
g1181 and n1435_not n1436_not ; n1437
g1182 and n1387_not n1437 ; n1438
g1183 and n1387 n1437_not ; n1439
g1184 and n1438_not n1439_not ; n1440
g1185 and n1386 n1440_not ; n1441
g1186 and n1386_not n1440 ; n1442
g1187 and n1441_not n1442_not ; n1443
g1188 and n1375_not n1443 ; n1444
g1189 and n1375 n1443_not ; n1445
g1190 and n1444_not n1445_not ; n1446
g1191 and n1374 n1446_not ; n1447
g1192 and n1374_not n1446 ; n1448
g1193 and n1447_not n1448_not ; n1449
g1194 and n1363_not n1449 ; n1450
g1195 and n1363 n1449_not ; n1451
g1196 and n1450_not n1451_not ; n1452
g1197 and n1362_not n1452 ; n1453
g1198 and n1452 n1453_not ; n1454
g1199 and n1362_not n1453_not ; n1455
g1200 and n1454_not n1455_not ; n1456
g1201 and n1243_not n1338 ; n1457
g1202 and n1342_not n1457_not ; n1458
g1203 and n1456_not n1458_not ; n1459
g1204 and n1456 n1458 ; n1460
g1205 and n1459_not n1460_not ; f[17]
g1206 and n1448_not n1450_not ; n1462
g1207 and b[15] n362 ; n1463
g1208 and b[13] n403 ; n1464
g1209 and b[14] n357 ; n1465
g1210 and n1464_not n1465_not ; n1466
g1211 and n1463_not n1466 ; n1467
g1212 and n365 n1131 ; n1468
g1213 and n1467 n1468_not ; n1469
g1214 and a[5] n1469_not ; n1470
g1215 and a[5] n1470_not ; n1471
g1216 and n1469_not n1470_not ; n1472
g1217 and n1471_not n1472_not ; n1473
g1218 and n1442_not n1444_not ; n1474
g1219 and b[12] n511 ; n1475
g1220 and b[10] n541 ; n1476
g1221 and b[11] n506 ; n1477
g1222 and n1476_not n1477_not ; n1478
g1223 and n1475_not n1478 ; n1479
g1224 and n514 n842 ; n1480
g1225 and n1479 n1480_not ; n1481
g1226 and a[8] n1481_not ; n1482
g1227 and a[8] n1482_not ; n1483
g1228 and n1481_not n1482_not ; n1484
g1229 and n1483_not n1484_not ; n1485
g1230 and n1436_not n1438_not ; n1486
g1231 and b[6] n951 ; n1487
g1232 and b[4] n1056 ; n1488
g1233 and b[5] n946 ; n1489
g1234 and n1488_not n1489_not ; n1490
g1235 and n1487_not n1490 ; n1491
g1236 and n459 n954 ; n1492
g1237 and n1491 n1492_not ; n1493
g1238 and a[14] n1493_not ; n1494
g1239 and a[14] n1494_not ; n1495
g1240 and n1493_not n1494_not ; n1496
g1241 and n1495_not n1496_not ; n1497
g1242 and a[17] a[18]_not ; n1498
g1243 and a[17]_not a[18] ; n1499
g1244 and n1498_not n1499_not ; n1500
g1245 and b[0] n1500_not ; n1501
g1246 and n1403_not n1501 ; n1502
g1247 and n1403 n1501_not ; n1503
g1248 and n1502_not n1503_not ; n1504
g1249 and b[3] n1302 ; n1505
g1250 and b[1] n1391 ; n1506
g1251 and b[2] n1297 ; n1507
g1252 and n1506_not n1507_not ; n1508
g1253 and n1505_not n1508 ; n1509
g1254 and n318 n1305 ; n1510
g1255 and n1509 n1510_not ; n1511
g1256 and a[17] n1511_not ; n1512
g1257 and a[17] n1512_not ; n1513
g1258 and n1511_not n1512_not ; n1514
g1259 and n1513_not n1514_not ; n1515
g1260 and n1504_not n1515_not ; n1516
g1261 and n1504 n1515 ; n1517
g1262 and n1516_not n1517_not ; n1518
g1263 and n1497_not n1518 ; n1519
g1264 and n1518 n1519_not ; n1520
g1265 and n1497_not n1519_not ; n1521
g1266 and n1520_not n1521_not ; n1522
g1267 and n1421_not n1522 ; n1523
g1268 and n1421 n1522_not ; n1524
g1269 and n1523_not n1524_not ; n1525
g1270 and b[9] n700 ; n1526
g1271 and b[7] n767 ; n1527
g1272 and b[8] n695 ; n1528
g1273 and n1527_not n1528_not ; n1529
g1274 and n1526_not n1529 ; n1530
g1275 and n651 n703 ; n1531
g1276 and n1530 n1531_not ; n1532
g1277 and a[11] n1532_not ; n1533
g1278 and a[11] n1533_not ; n1534
g1279 and n1532_not n1533_not ; n1535
g1280 and n1534_not n1535_not ; n1536
g1281 and n1525_not n1536_not ; n1537
g1282 and n1525 n1536 ; n1538
g1283 and n1537_not n1538_not ; n1539
g1284 and n1486_not n1539 ; n1540
g1285 and n1486 n1539_not ; n1541
g1286 and n1540_not n1541_not ; n1542
g1287 and n1485 n1542_not ; n1543
g1288 and n1485_not n1542 ; n1544
g1289 and n1543_not n1544_not ; n1545
g1290 and n1474_not n1545 ; n1546
g1291 and n1474 n1545_not ; n1547
g1292 and n1546_not n1547_not ; n1548
g1293 and n1473_not n1548 ; n1549
g1294 and n1473 n1548_not ; n1550
g1295 and n1549_not n1550_not ; n1551
g1296 and n1462_not n1551 ; n1552
g1297 and n1462 n1551_not ; n1553
g1298 and n1552_not n1553_not ; n1554
g1299 and b[18] n266 ; n1555
g1300 and b[16] n284 ; n1556
g1301 and b[17] n261 ; n1557
g1302 and n1556_not n1557_not ; n1558
g1303 and n1555_not n1558 ; n1559
g1304 and n1352_not n1354_not ; n1560
g1305 and b[17]_not b[18]_not ; n1561
g1306 and b[17] b[18] ; n1562
g1307 and n1561_not n1562_not ; n1563
g1308 and n1560_not n1563 ; n1564
g1309 and n1560 n1563_not ; n1565
g1310 and n1564_not n1565_not ; n1566
g1311 and n269 n1566 ; n1567
g1312 and n1559 n1567_not ; n1568
g1313 and a[2] n1568_not ; n1569
g1314 and a[2] n1569_not ; n1570
g1315 and n1568_not n1569_not ; n1571
g1316 and n1570_not n1571_not ; n1572
g1317 and n1554 n1572_not ; n1573
g1318 and n1554 n1573_not ; n1574
g1319 and n1572_not n1573_not ; n1575
g1320 and n1574_not n1575_not ; n1576
g1321 and n1453_not n1459_not ; n1577
g1322 and n1576_not n1577_not ; n1578
g1323 and n1576 n1577 ; n1579
g1324 and n1578_not n1579_not ; f[18]
g1325 and b[16] n362 ; n1581
g1326 and b[14] n403 ; n1582
g1327 and b[15] n357 ; n1583
g1328 and n1582_not n1583_not ; n1584
g1329 and n1581_not n1584 ; n1585
g1330 and n365 n1237 ; n1586
g1331 and n1585 n1586_not ; n1587
g1332 and a[5] n1587_not ; n1588
g1333 and a[5] n1588_not ; n1589
g1334 and n1587_not n1588_not ; n1590
g1335 and n1589_not n1590_not ; n1591
g1336 and n1421_not n1522_not ; n1592
g1337 and n1519_not n1592_not ; n1593
g1338 and b[7] n951 ; n1594
g1339 and b[5] n1056 ; n1595
g1340 and b[6] n946 ; n1596
g1341 and n1595_not n1596_not ; n1597
g1342 and n1594_not n1597 ; n1598
g1343 and n484 n954 ; n1599
g1344 and n1598 n1599_not ; n1600
g1345 and a[14] n1600_not ; n1601
g1346 and a[14] n1601_not ; n1602
g1347 and n1600_not n1601_not ; n1603
g1348 and n1602_not n1603_not ; n1604
g1349 and n1403 n1501 ; n1605
g1350 and n1516_not n1605_not ; n1606
g1351 and b[4] n1302 ; n1607
g1352 and b[2] n1391 ; n1608
g1353 and b[3] n1297 ; n1609
g1354 and n1608_not n1609_not ; n1610
g1355 and n1607_not n1610 ; n1611
g1356 and n346 n1305 ; n1612
g1357 and n1611 n1612_not ; n1613
g1358 and a[17] n1613_not ; n1614
g1359 and a[17] n1614_not ; n1615
g1360 and n1613_not n1614_not ; n1616
g1361 and n1615_not n1616_not ; n1617
g1362 and a[20] n1501_not ; n1618
g1363 and a[18]_not a[19] ; n1619
g1364 and a[18] a[19]_not ; n1620
g1365 and n1619_not n1620_not ; n1621
g1366 and n1500 n1621_not ; n1622
g1367 and b[0] n1622 ; n1623
g1368 and a[19]_not a[20] ; n1624
g1369 and a[19] a[20]_not ; n1625
g1370 and n1624_not n1625_not ; n1626
g1371 and n1500_not n1626 ; n1627
g1372 and b[1] n1627 ; n1628
g1373 and n1623_not n1628_not ; n1629
g1374 and n1500_not n1626_not ; n1630
g1375 and n272_not n1630 ; n1631
g1376 and n1629 n1631_not ; n1632
g1377 and a[20] n1632_not ; n1633
g1378 and a[20] n1633_not ; n1634
g1379 and n1632_not n1633_not ; n1635
g1380 and n1634_not n1635_not ; n1636
g1381 and n1618 n1636_not ; n1637
g1382 and n1618_not n1636 ; n1638
g1383 and n1637_not n1638_not ; n1639
g1384 and n1617 n1639 ; n1640
g1385 and n1617_not n1639_not ; n1641
g1386 and n1640_not n1641_not ; n1642
g1387 and n1606_not n1642_not ; n1643
g1388 and n1606 n1642 ; n1644
g1389 and n1643_not n1644_not ; n1645
g1390 and n1604_not n1645 ; n1646
g1391 and n1604 n1645_not ; n1647
g1392 and n1646_not n1647_not ; n1648
g1393 and n1593_not n1648 ; n1649
g1394 and n1593 n1648_not ; n1650
g1395 and n1649_not n1650_not ; n1651
g1396 and b[10] n700 ; n1652
g1397 and b[8] n767 ; n1653
g1398 and b[9] n695 ; n1654
g1399 and n1653_not n1654_not ; n1655
g1400 and n1652_not n1655 ; n1656
g1401 and n703 n738 ; n1657
g1402 and n1656 n1657_not ; n1658
g1403 and a[11] n1658_not ; n1659
g1404 and a[11] n1659_not ; n1660
g1405 and n1658_not n1659_not ; n1661
g1406 and n1660_not n1661_not ; n1662
g1407 and n1651 n1662_not ; n1663
g1408 and n1651 n1663_not ; n1664
g1409 and n1662_not n1663_not ; n1665
g1410 and n1664_not n1665_not ; n1666
g1411 and n1537_not n1540_not ; n1667
g1412 and n1666 n1667 ; n1668
g1413 and n1666_not n1667_not ; n1669
g1414 and n1668_not n1669_not ; n1670
g1415 and b[13] n511 ; n1671
g1416 and b[11] n541 ; n1672
g1417 and b[12] n506 ; n1673
g1418 and n1672_not n1673_not ; n1674
g1419 and n1671_not n1674 ; n1675
g1420 and n514 n1008 ; n1676
g1421 and n1675 n1676_not ; n1677
g1422 and a[8] n1677_not ; n1678
g1423 and a[8] n1678_not ; n1679
g1424 and n1677_not n1678_not ; n1680
g1425 and n1679_not n1680_not ; n1681
g1426 and n1670_not n1681 ; n1682
g1427 and n1670 n1681_not ; n1683
g1428 and n1682_not n1683_not ; n1684
g1429 and n1544_not n1546_not ; n1685
g1430 and n1684 n1685_not ; n1686
g1431 and n1684_not n1685 ; n1687
g1432 and n1686_not n1687_not ; n1688
g1433 and n1591_not n1688 ; n1689
g1434 and n1688 n1689_not ; n1690
g1435 and n1591_not n1689_not ; n1691
g1436 and n1690_not n1691_not ; n1692
g1437 and n1549_not n1552_not ; n1693
g1438 and n1692 n1693 ; n1694
g1439 and n1692_not n1693_not ; n1695
g1440 and n1694_not n1695_not ; n1696
g1441 and b[19] n266 ; n1697
g1442 and b[17] n284 ; n1698
g1443 and b[18] n261 ; n1699
g1444 and n1698_not n1699_not ; n1700
g1445 and n1697_not n1700 ; n1701
g1446 and n1562_not n1564_not ; n1702
g1447 and b[18]_not b[19]_not ; n1703
g1448 and b[18] b[19] ; n1704
g1449 and n1703_not n1704_not ; n1705
g1450 and n1702_not n1705 ; n1706
g1451 and n1702 n1705_not ; n1707
g1452 and n1706_not n1707_not ; n1708
g1453 and n269 n1708 ; n1709
g1454 and n1701 n1709_not ; n1710
g1455 and a[2] n1710_not ; n1711
g1456 and a[2] n1711_not ; n1712
g1457 and n1710_not n1711_not ; n1713
g1458 and n1712_not n1713_not ; n1714
g1459 and n1696 n1714_not ; n1715
g1460 and n1696 n1715_not ; n1716
g1461 and n1714_not n1715_not ; n1717
g1462 and n1716_not n1717_not ; n1718
g1463 and n1573_not n1578_not ; n1719
g1464 and n1718_not n1719_not ; n1720
g1465 and n1718 n1719 ; n1721
g1466 and n1720_not n1721_not ; f[19]
g1467 and n1689_not n1695_not ; n1723
g1468 and b[17] n362 ; n1724
g1469 and b[15] n403 ; n1725
g1470 and b[16] n357 ; n1726
g1471 and n1725_not n1726_not ; n1727
g1472 and n1724_not n1727 ; n1728
g1473 and n365 n1356 ; n1729
g1474 and n1728 n1729_not ; n1730
g1475 and a[5] n1730_not ; n1731
g1476 and a[5] n1731_not ; n1732
g1477 and n1730_not n1731_not ; n1733
g1478 and n1732_not n1733_not ; n1734
g1479 and b[14] n511 ; n1735
g1480 and b[12] n541 ; n1736
g1481 and b[13] n506 ; n1737
g1482 and n1736_not n1737_not ; n1738
g1483 and n1735_not n1738 ; n1739
g1484 and n514 n1034 ; n1740
g1485 and n1739 n1740_not ; n1741
g1486 and a[8] n1741_not ; n1742
g1487 and a[8] n1742_not ; n1743
g1488 and n1741_not n1742_not ; n1744
g1489 and n1743_not n1744_not ; n1745
g1490 and n1663_not n1669_not ; n1746
g1491 and b[11] n700 ; n1747
g1492 and b[9] n767 ; n1748
g1493 and b[10] n695 ; n1749
g1494 and n1748_not n1749_not ; n1750
g1495 and n1747_not n1750 ; n1751
g1496 and n703 n818 ; n1752
g1497 and n1751 n1752_not ; n1753
g1498 and a[11] n1753_not ; n1754
g1499 and a[11] n1754_not ; n1755
g1500 and n1753_not n1754_not ; n1756
g1501 and n1755_not n1756_not ; n1757
g1502 and n1646_not n1649_not ; n1758
g1503 and n1617_not n1639 ; n1759
g1504 and n1643_not n1759_not ; n1760
g1505 and b[2] n1627 ; n1761
g1506 and n1500 n1626_not ; n1762
g1507 and n1621 n1762 ; n1763
g1508 and b[0] n1763 ; n1764
g1509 and b[1] n1622 ; n1765
g1510 and n1764_not n1765_not ; n1766
g1511 and n1761_not n1766 ; n1767
g1512 and n296 n1630 ; n1768
g1513 and n1767 n1768_not ; n1769
g1514 and a[20] n1769_not ; n1770
g1515 and a[20] n1770_not ; n1771
g1516 and n1769_not n1770_not ; n1772
g1517 and n1771_not n1772_not ; n1773
g1518 and n1637_not n1773 ; n1774
g1519 and n1637 n1773_not ; n1775
g1520 and n1774_not n1775_not ; n1776
g1521 and b[5] n1302 ; n1777
g1522 and b[3] n1391 ; n1778
g1523 and b[4] n1297 ; n1779
g1524 and n1778_not n1779_not ; n1780
g1525 and n1777_not n1780 ; n1781
g1526 and n394 n1305 ; n1782
g1527 and n1781 n1782_not ; n1783
g1528 and a[17] n1783_not ; n1784
g1529 and a[17] n1784_not ; n1785
g1530 and n1783_not n1784_not ; n1786
g1531 and n1785_not n1786_not ; n1787
g1532 and n1776 n1787_not ; n1788
g1533 and n1776_not n1787 ; n1789
g1534 and n1760_not n1789_not ; n1790
g1535 and n1788_not n1790 ; n1791
g1536 and n1760_not n1791_not ; n1792
g1537 and n1788_not n1791_not ; n1793
g1538 and n1789_not n1793 ; n1794
g1539 and n1792_not n1794_not ; n1795
g1540 and b[8] n951 ; n1796
g1541 and b[6] n1056 ; n1797
g1542 and b[7] n946 ; n1798
g1543 and n1797_not n1798_not ; n1799
g1544 and n1796_not n1799 ; n1800
g1545 and n585 n954 ; n1801
g1546 and n1800 n1801_not ; n1802
g1547 and a[14] n1802_not ; n1803
g1548 and a[14] n1803_not ; n1804
g1549 and n1802_not n1803_not ; n1805
g1550 and n1804_not n1805_not ; n1806
g1551 and n1795 n1806 ; n1807
g1552 and n1795_not n1806_not ; n1808
g1553 and n1807_not n1808_not ; n1809
g1554 and n1758_not n1809 ; n1810
g1555 and n1758 n1809_not ; n1811
g1556 and n1810_not n1811_not ; n1812
g1557 and n1757 n1812_not ; n1813
g1558 and n1757_not n1812 ; n1814
g1559 and n1813_not n1814_not ; n1815
g1560 and n1746_not n1815 ; n1816
g1561 and n1746 n1815_not ; n1817
g1562 and n1816_not n1817_not ; n1818
g1563 and n1745_not n1818 ; n1819
g1564 and n1818 n1819_not ; n1820
g1565 and n1745_not n1819_not ; n1821
g1566 and n1820_not n1821_not ; n1822
g1567 and n1683_not n1686_not ; n1823
g1568 and n1822_not n1823_not ; n1824
g1569 and n1822 n1823 ; n1825
g1570 and n1824_not n1825_not ; n1826
g1571 and n1734_not n1826 ; n1827
g1572 and n1734_not n1827_not ; n1828
g1573 and n1826 n1827_not ; n1829
g1574 and n1828_not n1829_not ; n1830
g1575 and n1723_not n1830_not ; n1831
g1576 and n1723_not n1831_not ; n1832
g1577 and n1830_not n1831_not ; n1833
g1578 and n1832_not n1833_not ; n1834
g1579 and b[20] n266 ; n1835
g1580 and b[18] n284 ; n1836
g1581 and b[19] n261 ; n1837
g1582 and n1836_not n1837_not ; n1838
g1583 and n1835_not n1838 ; n1839
g1584 and n1704_not n1706_not ; n1840
g1585 and b[19]_not b[20]_not ; n1841
g1586 and b[19] b[20] ; n1842
g1587 and n1841_not n1842_not ; n1843
g1588 and n1840_not n1843 ; n1844
g1589 and n1840 n1843_not ; n1845
g1590 and n1844_not n1845_not ; n1846
g1591 and n269 n1846 ; n1847
g1592 and n1839 n1847_not ; n1848
g1593 and a[2] n1848_not ; n1849
g1594 and a[2] n1849_not ; n1850
g1595 and n1848_not n1849_not ; n1851
g1596 and n1850_not n1851_not ; n1852
g1597 and n1834_not n1852_not ; n1853
g1598 and n1834_not n1853_not ; n1854
g1599 and n1852_not n1853_not ; n1855
g1600 and n1854_not n1855_not ; n1856
g1601 and n1715_not n1720_not ; n1857
g1602 and n1856_not n1857_not ; n1858
g1603 and n1856 n1857 ; n1859
g1604 and n1858_not n1859_not ; f[20]
g1605 and n1819_not n1824_not ; n1861
g1606 and b[15] n511 ; n1862
g1607 and b[13] n541 ; n1863
g1608 and b[14] n506 ; n1864
g1609 and n1863_not n1864_not ; n1865
g1610 and n1862_not n1865 ; n1866
g1611 and n514 n1131 ; n1867
g1612 and n1866 n1867_not ; n1868
g1613 and a[8] n1868_not ; n1869
g1614 and a[8] n1869_not ; n1870
g1615 and n1868_not n1869_not ; n1871
g1616 and n1870_not n1871_not ; n1872
g1617 and n1814_not n1816_not ; n1873
g1618 and b[12] n700 ; n1874
g1619 and b[10] n767 ; n1875
g1620 and b[11] n695 ; n1876
g1621 and n1875_not n1876_not ; n1877
g1622 and n1874_not n1877 ; n1878
g1623 and n703 n842 ; n1879
g1624 and n1878 n1879_not ; n1880
g1625 and a[11] n1880_not ; n1881
g1626 and a[11] n1881_not ; n1882
g1627 and n1880_not n1881_not ; n1883
g1628 and n1882_not n1883_not ; n1884
g1629 and n1808_not n1810_not ; n1885
g1630 and b[6] n1302 ; n1886
g1631 and b[4] n1391 ; n1887
g1632 and b[5] n1297 ; n1888
g1633 and n1887_not n1888_not ; n1889
g1634 and n1886_not n1889 ; n1890
g1635 and n459 n1305 ; n1891
g1636 and n1890 n1891_not ; n1892
g1637 and a[17] n1892_not ; n1893
g1638 and a[17] n1893_not ; n1894
g1639 and n1892_not n1893_not ; n1895
g1640 and n1894_not n1895_not ; n1896
g1641 and a[20] a[21]_not ; n1897
g1642 and a[20]_not a[21] ; n1898
g1643 and n1897_not n1898_not ; n1899
g1644 and b[0] n1899_not ; n1900
g1645 and n1775_not n1900 ; n1901
g1646 and n1775 n1900_not ; n1902
g1647 and n1901_not n1902_not ; n1903
g1648 and b[3] n1627 ; n1904
g1649 and b[1] n1763 ; n1905
g1650 and b[2] n1622 ; n1906
g1651 and n1905_not n1906_not ; n1907
g1652 and n1904_not n1907 ; n1908
g1653 and n318 n1630 ; n1909
g1654 and n1908 n1909_not ; n1910
g1655 and a[20] n1910_not ; n1911
g1656 and a[20] n1911_not ; n1912
g1657 and n1910_not n1911_not ; n1913
g1658 and n1912_not n1913_not ; n1914
g1659 and n1903_not n1914_not ; n1915
g1660 and n1903 n1914 ; n1916
g1661 and n1915_not n1916_not ; n1917
g1662 and n1896_not n1917 ; n1918
g1663 and n1917 n1918_not ; n1919
g1664 and n1896_not n1918_not ; n1920
g1665 and n1919_not n1920_not ; n1921
g1666 and n1793_not n1921 ; n1922
g1667 and n1793 n1921_not ; n1923
g1668 and n1922_not n1923_not ; n1924
g1669 and b[9] n951 ; n1925
g1670 and b[7] n1056 ; n1926
g1671 and b[8] n946 ; n1927
g1672 and n1926_not n1927_not ; n1928
g1673 and n1925_not n1928 ; n1929
g1674 and n651 n954 ; n1930
g1675 and n1929 n1930_not ; n1931
g1676 and a[14] n1931_not ; n1932
g1677 and a[14] n1932_not ; n1933
g1678 and n1931_not n1932_not ; n1934
g1679 and n1933_not n1934_not ; n1935
g1680 and n1924_not n1935_not ; n1936
g1681 and n1924 n1935 ; n1937
g1682 and n1936_not n1937_not ; n1938
g1683 and n1885_not n1938 ; n1939
g1684 and n1885 n1938_not ; n1940
g1685 and n1939_not n1940_not ; n1941
g1686 and n1884 n1941_not ; n1942
g1687 and n1884_not n1941 ; n1943
g1688 and n1942_not n1943_not ; n1944
g1689 and n1873_not n1944 ; n1945
g1690 and n1873 n1944_not ; n1946
g1691 and n1945_not n1946_not ; n1947
g1692 and n1872_not n1947 ; n1948
g1693 and n1872 n1947_not ; n1949
g1694 and n1948_not n1949_not ; n1950
g1695 and n1861_not n1950 ; n1951
g1696 and n1861 n1950_not ; n1952
g1697 and n1951_not n1952_not ; n1953
g1698 and b[18] n362 ; n1954
g1699 and b[16] n403 ; n1955
g1700 and b[17] n357 ; n1956
g1701 and n1955_not n1956_not ; n1957
g1702 and n1954_not n1957 ; n1958
g1703 and n365 n1566 ; n1959
g1704 and n1958 n1959_not ; n1960
g1705 and a[5] n1960_not ; n1961
g1706 and a[5] n1961_not ; n1962
g1707 and n1960_not n1961_not ; n1963
g1708 and n1962_not n1963_not ; n1964
g1709 and n1953 n1964_not ; n1965
g1710 and n1953 n1965_not ; n1966
g1711 and n1964_not n1965_not ; n1967
g1712 and n1966_not n1967_not ; n1968
g1713 and n1827_not n1831_not ; n1969
g1714 and n1968 n1969 ; n1970
g1715 and n1968_not n1969_not ; n1971
g1716 and n1970_not n1971_not ; n1972
g1717 and b[21] n266 ; n1973
g1718 and b[19] n284 ; n1974
g1719 and b[20] n261 ; n1975
g1720 and n1974_not n1975_not ; n1976
g1721 and n1973_not n1976 ; n1977
g1722 and n1842_not n1844_not ; n1978
g1723 and b[20]_not b[21]_not ; n1979
g1724 and b[20] b[21] ; n1980
g1725 and n1979_not n1980_not ; n1981
g1726 and n1978_not n1981 ; n1982
g1727 and n1978 n1981_not ; n1983
g1728 and n1982_not n1983_not ; n1984
g1729 and n269 n1984 ; n1985
g1730 and n1977 n1985_not ; n1986
g1731 and a[2] n1986_not ; n1987
g1732 and a[2] n1987_not ; n1988
g1733 and n1986_not n1987_not ; n1989
g1734 and n1988_not n1989_not ; n1990
g1735 and n1972 n1990_not ; n1991
g1736 and n1972 n1991_not ; n1992
g1737 and n1990_not n1991_not ; n1993
g1738 and n1992_not n1993_not ; n1994
g1739 and n1853_not n1858_not ; n1995
g1740 and n1994_not n1995_not ; n1996
g1741 and n1994 n1995 ; n1997
g1742 and n1996_not n1997_not ; f[21]
g1743 and n1991_not n1996_not ; n1999
g1744 and n1948_not n1951_not ; n2000
g1745 and b[16] n511 ; n2001
g1746 and b[14] n541 ; n2002
g1747 and b[15] n506 ; n2003
g1748 and n2002_not n2003_not ; n2004
g1749 and n2001_not n2004 ; n2005
g1750 and n514 n1237 ; n2006
g1751 and n2005 n2006_not ; n2007
g1752 and a[8] n2007_not ; n2008
g1753 and a[8] n2008_not ; n2009
g1754 and n2007_not n2008_not ; n2010
g1755 and n2009_not n2010_not ; n2011
g1756 and n1943_not n1945_not ; n2012
g1757 and n1793_not n1921_not ; n2013
g1758 and n1918_not n2013_not ; n2014
g1759 and b[7] n1302 ; n2015
g1760 and b[5] n1391 ; n2016
g1761 and b[6] n1297 ; n2017
g1762 and n2016_not n2017_not ; n2018
g1763 and n2015_not n2018 ; n2019
g1764 and n484 n1305 ; n2020
g1765 and n2019 n2020_not ; n2021
g1766 and a[17] n2021_not ; n2022
g1767 and a[17] n2022_not ; n2023
g1768 and n2021_not n2022_not ; n2024
g1769 and n2023_not n2024_not ; n2025
g1770 and n1775 n1900 ; n2026
g1771 and n1915_not n2026_not ; n2027
g1772 and b[4] n1627 ; n2028
g1773 and b[2] n1763 ; n2029
g1774 and b[3] n1622 ; n2030
g1775 and n2029_not n2030_not ; n2031
g1776 and n2028_not n2031 ; n2032
g1777 and n346 n1630 ; n2033
g1778 and n2032 n2033_not ; n2034
g1779 and a[20] n2034_not ; n2035
g1780 and a[20] n2035_not ; n2036
g1781 and n2034_not n2035_not ; n2037
g1782 and n2036_not n2037_not ; n2038
g1783 and a[23] n1900_not ; n2039
g1784 and a[21]_not a[22] ; n2040
g1785 and a[21] a[22]_not ; n2041
g1786 and n2040_not n2041_not ; n2042
g1787 and n1899 n2042_not ; n2043
g1788 and b[0] n2043 ; n2044
g1789 and a[22]_not a[23] ; n2045
g1790 and a[22] a[23]_not ; n2046
g1791 and n2045_not n2046_not ; n2047
g1792 and n1899_not n2047 ; n2048
g1793 and b[1] n2048 ; n2049
g1794 and n2044_not n2049_not ; n2050
g1795 and n1899_not n2047_not ; n2051
g1796 and n272_not n2051 ; n2052
g1797 and n2050 n2052_not ; n2053
g1798 and a[23] n2053_not ; n2054
g1799 and a[23] n2054_not ; n2055
g1800 and n2053_not n2054_not ; n2056
g1801 and n2055_not n2056_not ; n2057
g1802 and n2039 n2057_not ; n2058
g1803 and n2039_not n2057 ; n2059
g1804 and n2058_not n2059_not ; n2060
g1805 and n2038 n2060 ; n2061
g1806 and n2038_not n2060_not ; n2062
g1807 and n2061_not n2062_not ; n2063
g1808 and n2027_not n2063_not ; n2064
g1809 and n2027 n2063 ; n2065
g1810 and n2064_not n2065_not ; n2066
g1811 and n2025_not n2066 ; n2067
g1812 and n2025 n2066_not ; n2068
g1813 and n2067_not n2068_not ; n2069
g1814 and n2014_not n2069 ; n2070
g1815 and n2014 n2069_not ; n2071
g1816 and n2070_not n2071_not ; n2072
g1817 and b[10] n951 ; n2073
g1818 and b[8] n1056 ; n2074
g1819 and b[9] n946 ; n2075
g1820 and n2074_not n2075_not ; n2076
g1821 and n2073_not n2076 ; n2077
g1822 and n738 n954 ; n2078
g1823 and n2077 n2078_not ; n2079
g1824 and a[14] n2079_not ; n2080
g1825 and a[14] n2080_not ; n2081
g1826 and n2079_not n2080_not ; n2082
g1827 and n2081_not n2082_not ; n2083
g1828 and n2072 n2083_not ; n2084
g1829 and n2072 n2084_not ; n2085
g1830 and n2083_not n2084_not ; n2086
g1831 and n2085_not n2086_not ; n2087
g1832 and n1936_not n1939_not ; n2088
g1833 and n2087 n2088 ; n2089
g1834 and n2087_not n2088_not ; n2090
g1835 and n2089_not n2090_not ; n2091
g1836 and b[13] n700 ; n2092
g1837 and b[11] n767 ; n2093
g1838 and b[12] n695 ; n2094
g1839 and n2093_not n2094_not ; n2095
g1840 and n2092_not n2095 ; n2096
g1841 and n703 n1008 ; n2097
g1842 and n2096 n2097_not ; n2098
g1843 and a[11] n2098_not ; n2099
g1844 and a[11] n2099_not ; n2100
g1845 and n2098_not n2099_not ; n2101
g1846 and n2100_not n2101_not ; n2102
g1847 and n2091_not n2102 ; n2103
g1848 and n2091 n2102_not ; n2104
g1849 and n2103_not n2104_not ; n2105
g1850 and n2012_not n2105 ; n2106
g1851 and n2012 n2105_not ; n2107
g1852 and n2106_not n2107_not ; n2108
g1853 and n2011_not n2108 ; n2109
g1854 and n2011 n2108_not ; n2110
g1855 and n2109_not n2110_not ; n2111
g1856 and n2000_not n2111 ; n2112
g1857 and n2000 n2111_not ; n2113
g1858 and n2112_not n2113_not ; n2114
g1859 and b[19] n362 ; n2115
g1860 and b[17] n403 ; n2116
g1861 and b[18] n357 ; n2117
g1862 and n2116_not n2117_not ; n2118
g1863 and n2115_not n2118 ; n2119
g1864 and n365 n1708 ; n2120
g1865 and n2119 n2120_not ; n2121
g1866 and a[5] n2121_not ; n2122
g1867 and a[5] n2122_not ; n2123
g1868 and n2121_not n2122_not ; n2124
g1869 and n2123_not n2124_not ; n2125
g1870 and n2114 n2125_not ; n2126
g1871 and n2114 n2126_not ; n2127
g1872 and n2125_not n2126_not ; n2128
g1873 and n2127_not n2128_not ; n2129
g1874 and n1965_not n1971_not ; n2130
g1875 and n2129 n2130 ; n2131
g1876 and n2129_not n2130_not ; n2132
g1877 and n2131_not n2132_not ; n2133
g1878 and b[22] n266 ; n2134
g1879 and b[20] n284 ; n2135
g1880 and b[21] n261 ; n2136
g1881 and n2135_not n2136_not ; n2137
g1882 and n2134_not n2137 ; n2138
g1883 and n1980_not n1982_not ; n2139
g1884 and b[21]_not b[22]_not ; n2140
g1885 and b[21] b[22] ; n2141
g1886 and n2140_not n2141_not ; n2142
g1887 and n2139_not n2142 ; n2143
g1888 and n2139 n2142_not ; n2144
g1889 and n2143_not n2144_not ; n2145
g1890 and n269 n2145 ; n2146
g1891 and n2138 n2146_not ; n2147
g1892 and a[2] n2147_not ; n2148
g1893 and a[2] n2148_not ; n2149
g1894 and n2147_not n2148_not ; n2150
g1895 and n2149_not n2150_not ; n2151
g1896 and n2133_not n2151 ; n2152
g1897 and n2133 n2151_not ; n2153
g1898 and n2152_not n2153_not ; n2154
g1899 and n1999_not n2154 ; n2155
g1900 and n1999 n2154_not ; n2156
g1901 and n2155_not n2156_not ; f[22]
g1902 and n2109_not n2112_not ; n2158
g1903 and b[17] n511 ; n2159
g1904 and b[15] n541 ; n2160
g1905 and b[16] n506 ; n2161
g1906 and n2160_not n2161_not ; n2162
g1907 and n2159_not n2162 ; n2163
g1908 and n514 n1356 ; n2164
g1909 and n2163 n2164_not ; n2165
g1910 and a[8] n2165_not ; n2166
g1911 and a[8] n2166_not ; n2167
g1912 and n2165_not n2166_not ; n2168
g1913 and n2167_not n2168_not ; n2169
g1914 and b[14] n700 ; n2170
g1915 and b[12] n767 ; n2171
g1916 and b[13] n695 ; n2172
g1917 and n2171_not n2172_not ; n2173
g1918 and n2170_not n2173 ; n2174
g1919 and n703 n1034 ; n2175
g1920 and n2174 n2175_not ; n2176
g1921 and a[11] n2176_not ; n2177
g1922 and a[11] n2177_not ; n2178
g1923 and n2176_not n2177_not ; n2179
g1924 and n2178_not n2179_not ; n2180
g1925 and n2084_not n2090_not ; n2181
g1926 and b[11] n951 ; n2182
g1927 and b[9] n1056 ; n2183
g1928 and b[10] n946 ; n2184
g1929 and n2183_not n2184_not ; n2185
g1930 and n2182_not n2185 ; n2186
g1931 and n818 n954 ; n2187
g1932 and n2186 n2187_not ; n2188
g1933 and a[14] n2188_not ; n2189
g1934 and a[14] n2189_not ; n2190
g1935 and n2188_not n2189_not ; n2191
g1936 and n2190_not n2191_not ; n2192
g1937 and n2067_not n2070_not ; n2193
g1938 and n2038_not n2060 ; n2194
g1939 and n2064_not n2194_not ; n2195
g1940 and b[2] n2048 ; n2196
g1941 and n1899 n2047_not ; n2197
g1942 and n2042 n2197 ; n2198
g1943 and b[0] n2198 ; n2199
g1944 and b[1] n2043 ; n2200
g1945 and n2199_not n2200_not ; n2201
g1946 and n2196_not n2201 ; n2202
g1947 and n296 n2051 ; n2203
g1948 and n2202 n2203_not ; n2204
g1949 and a[23] n2204_not ; n2205
g1950 and a[23] n2205_not ; n2206
g1951 and n2204_not n2205_not ; n2207
g1952 and n2206_not n2207_not ; n2208
g1953 and n2058_not n2208 ; n2209
g1954 and n2058 n2208_not ; n2210
g1955 and n2209_not n2210_not ; n2211
g1956 and b[5] n1627 ; n2212
g1957 and b[3] n1763 ; n2213
g1958 and b[4] n1622 ; n2214
g1959 and n2213_not n2214_not ; n2215
g1960 and n2212_not n2215 ; n2216
g1961 and n394 n1630 ; n2217
g1962 and n2216 n2217_not ; n2218
g1963 and a[20] n2218_not ; n2219
g1964 and a[20] n2219_not ; n2220
g1965 and n2218_not n2219_not ; n2221
g1966 and n2220_not n2221_not ; n2222
g1967 and n2211 n2222_not ; n2223
g1968 and n2211_not n2222 ; n2224
g1969 and n2195_not n2224_not ; n2225
g1970 and n2223_not n2225 ; n2226
g1971 and n2195_not n2226_not ; n2227
g1972 and n2223_not n2226_not ; n2228
g1973 and n2224_not n2228 ; n2229
g1974 and n2227_not n2229_not ; n2230
g1975 and b[8] n1302 ; n2231
g1976 and b[6] n1391 ; n2232
g1977 and b[7] n1297 ; n2233
g1978 and n2232_not n2233_not ; n2234
g1979 and n2231_not n2234 ; n2235
g1980 and n585 n1305 ; n2236
g1981 and n2235 n2236_not ; n2237
g1982 and a[17] n2237_not ; n2238
g1983 and a[17] n2238_not ; n2239
g1984 and n2237_not n2238_not ; n2240
g1985 and n2239_not n2240_not ; n2241
g1986 and n2230 n2241 ; n2242
g1987 and n2230_not n2241_not ; n2243
g1988 and n2242_not n2243_not ; n2244
g1989 and n2193_not n2244 ; n2245
g1990 and n2193 n2244_not ; n2246
g1991 and n2245_not n2246_not ; n2247
g1992 and n2192 n2247_not ; n2248
g1993 and n2192_not n2247 ; n2249
g1994 and n2248_not n2249_not ; n2250
g1995 and n2181_not n2250 ; n2251
g1996 and n2181 n2250_not ; n2252
g1997 and n2251_not n2252_not ; n2253
g1998 and n2180_not n2253 ; n2254
g1999 and n2253 n2254_not ; n2255
g2000 and n2180_not n2254_not ; n2256
g2001 and n2255_not n2256_not ; n2257
g2002 and n2104_not n2106_not ; n2258
g2003 and n2257_not n2258_not ; n2259
g2004 and n2257 n2258 ; n2260
g2005 and n2259_not n2260_not ; n2261
g2006 and n2169_not n2261 ; n2262
g2007 and n2169_not n2262_not ; n2263
g2008 and n2261 n2262_not ; n2264
g2009 and n2263_not n2264_not ; n2265
g2010 and n2158_not n2265_not ; n2266
g2011 and n2158_not n2266_not ; n2267
g2012 and n2265_not n2266_not ; n2268
g2013 and n2267_not n2268_not ; n2269
g2014 and b[20] n362 ; n2270
g2015 and b[18] n403 ; n2271
g2016 and b[19] n357 ; n2272
g2017 and n2271_not n2272_not ; n2273
g2018 and n2270_not n2273 ; n2274
g2019 and n365 n1846 ; n2275
g2020 and n2274 n2275_not ; n2276
g2021 and a[5] n2276_not ; n2277
g2022 and a[5] n2277_not ; n2278
g2023 and n2276_not n2277_not ; n2279
g2024 and n2278_not n2279_not ; n2280
g2025 and n2269_not n2280_not ; n2281
g2026 and n2269_not n2281_not ; n2282
g2027 and n2280_not n2281_not ; n2283
g2028 and n2282_not n2283_not ; n2284
g2029 and n2126_not n2132_not ; n2285
g2030 and n2284 n2285 ; n2286
g2031 and n2284_not n2285_not ; n2287
g2032 and n2286_not n2287_not ; n2288
g2033 and b[23] n266 ; n2289
g2034 and b[21] n284 ; n2290
g2035 and b[22] n261 ; n2291
g2036 and n2290_not n2291_not ; n2292
g2037 and n2289_not n2292 ; n2293
g2038 and n2141_not n2143_not ; n2294
g2039 and b[22]_not b[23]_not ; n2295
g2040 and b[22] b[23] ; n2296
g2041 and n2295_not n2296_not ; n2297
g2042 and n2294_not n2297 ; n2298
g2043 and n2294 n2297_not ; n2299
g2044 and n2298_not n2299_not ; n2300
g2045 and n269 n2300 ; n2301
g2046 and n2293 n2301_not ; n2302
g2047 and a[2] n2302_not ; n2303
g2048 and a[2] n2303_not ; n2304
g2049 and n2302_not n2303_not ; n2305
g2050 and n2304_not n2305_not ; n2306
g2051 and n2288 n2306_not ; n2307
g2052 and n2288 n2307_not ; n2308
g2053 and n2306_not n2307_not ; n2309
g2054 and n2308_not n2309_not ; n2310
g2055 and n2153_not n2155_not ; n2311
g2056 and n2310_not n2311_not ; n2312
g2057 and n2310 n2311 ; n2313
g2058 and n2312_not n2313_not ; f[23]
g2059 and n2281_not n2287_not ; n2315
g2060 and b[21] n362 ; n2316
g2061 and b[19] n403 ; n2317
g2062 and b[20] n357 ; n2318
g2063 and n2317_not n2318_not ; n2319
g2064 and n2316_not n2319 ; n2320
g2065 and n365 n1984 ; n2321
g2066 and n2320 n2321_not ; n2322
g2067 and a[5] n2322_not ; n2323
g2068 and a[5] n2323_not ; n2324
g2069 and n2322_not n2323_not ; n2325
g2070 and n2324_not n2325_not ; n2326
g2071 and n2262_not n2266_not ; n2327
g2072 and b[15] n700 ; n2328
g2073 and b[13] n767 ; n2329
g2074 and b[14] n695 ; n2330
g2075 and n2329_not n2330_not ; n2331
g2076 and n2328_not n2331 ; n2332
g2077 and n703 n1131 ; n2333
g2078 and n2332 n2333_not ; n2334
g2079 and a[11] n2334_not ; n2335
g2080 and a[11] n2335_not ; n2336
g2081 and n2334_not n2335_not ; n2337
g2082 and n2336_not n2337_not ; n2338
g2083 and n2249_not n2251_not ; n2339
g2084 and b[12] n951 ; n2340
g2085 and b[10] n1056 ; n2341
g2086 and b[11] n946 ; n2342
g2087 and n2341_not n2342_not ; n2343
g2088 and n2340_not n2343 ; n2344
g2089 and n842 n954 ; n2345
g2090 and n2344 n2345_not ; n2346
g2091 and a[14] n2346_not ; n2347
g2092 and a[14] n2347_not ; n2348
g2093 and n2346_not n2347_not ; n2349
g2094 and n2348_not n2349_not ; n2350
g2095 and n2243_not n2245_not ; n2351
g2096 and b[6] n1627 ; n2352
g2097 and b[4] n1763 ; n2353
g2098 and b[5] n1622 ; n2354
g2099 and n2353_not n2354_not ; n2355
g2100 and n2352_not n2355 ; n2356
g2101 and n459 n1630 ; n2357
g2102 and n2356 n2357_not ; n2358
g2103 and a[20] n2358_not ; n2359
g2104 and a[20] n2359_not ; n2360
g2105 and n2358_not n2359_not ; n2361
g2106 and n2360_not n2361_not ; n2362
g2107 and a[23] a[24]_not ; n2363
g2108 and a[23]_not a[24] ; n2364
g2109 and n2363_not n2364_not ; n2365
g2110 and b[0] n2365_not ; n2366
g2111 and n2210_not n2366 ; n2367
g2112 and n2210 n2366_not ; n2368
g2113 and n2367_not n2368_not ; n2369
g2114 and b[3] n2048 ; n2370
g2115 and b[1] n2198 ; n2371
g2116 and b[2] n2043 ; n2372
g2117 and n2371_not n2372_not ; n2373
g2118 and n2370_not n2373 ; n2374
g2119 and n318 n2051 ; n2375
g2120 and n2374 n2375_not ; n2376
g2121 and a[23] n2376_not ; n2377
g2122 and a[23] n2377_not ; n2378
g2123 and n2376_not n2377_not ; n2379
g2124 and n2378_not n2379_not ; n2380
g2125 and n2369_not n2380_not ; n2381
g2126 and n2369 n2380 ; n2382
g2127 and n2381_not n2382_not ; n2383
g2128 and n2362_not n2383 ; n2384
g2129 and n2383 n2384_not ; n2385
g2130 and n2362_not n2384_not ; n2386
g2131 and n2385_not n2386_not ; n2387
g2132 and n2228_not n2387 ; n2388
g2133 and n2228 n2387_not ; n2389
g2134 and n2388_not n2389_not ; n2390
g2135 and b[9] n1302 ; n2391
g2136 and b[7] n1391 ; n2392
g2137 and b[8] n1297 ; n2393
g2138 and n2392_not n2393_not ; n2394
g2139 and n2391_not n2394 ; n2395
g2140 and n651 n1305 ; n2396
g2141 and n2395 n2396_not ; n2397
g2142 and a[17] n2397_not ; n2398
g2143 and a[17] n2398_not ; n2399
g2144 and n2397_not n2398_not ; n2400
g2145 and n2399_not n2400_not ; n2401
g2146 and n2390_not n2401_not ; n2402
g2147 and n2390 n2401 ; n2403
g2148 and n2402_not n2403_not ; n2404
g2149 and n2351_not n2404 ; n2405
g2150 and n2351 n2404_not ; n2406
g2151 and n2405_not n2406_not ; n2407
g2152 and n2350 n2407_not ; n2408
g2153 and n2350_not n2407 ; n2409
g2154 and n2408_not n2409_not ; n2410
g2155 and n2339_not n2410 ; n2411
g2156 and n2339 n2410_not ; n2412
g2157 and n2411_not n2412_not ; n2413
g2158 and n2338_not n2413 ; n2414
g2159 and n2413 n2414_not ; n2415
g2160 and n2338_not n2414_not ; n2416
g2161 and n2415_not n2416_not ; n2417
g2162 and n2254_not n2259_not ; n2418
g2163 and n2417 n2418 ; n2419
g2164 and n2417_not n2418_not ; n2420
g2165 and n2419_not n2420_not ; n2421
g2166 and b[18] n511 ; n2422
g2167 and b[16] n541 ; n2423
g2168 and b[17] n506 ; n2424
g2169 and n2423_not n2424_not ; n2425
g2170 and n2422_not n2425 ; n2426
g2171 and n514 n1566 ; n2427
g2172 and n2426 n2427_not ; n2428
g2173 and a[8] n2428_not ; n2429
g2174 and a[8] n2429_not ; n2430
g2175 and n2428_not n2429_not ; n2431
g2176 and n2430_not n2431_not ; n2432
g2177 and n2421_not n2432 ; n2433
g2178 and n2421 n2432_not ; n2434
g2179 and n2433_not n2434_not ; n2435
g2180 and n2327_not n2435 ; n2436
g2181 and n2327 n2435_not ; n2437
g2182 and n2436_not n2437_not ; n2438
g2183 and n2326_not n2438 ; n2439
g2184 and n2326_not n2439_not ; n2440
g2185 and n2438 n2439_not ; n2441
g2186 and n2440_not n2441_not ; n2442
g2187 and n2315_not n2442_not ; n2443
g2188 and n2315_not n2443_not ; n2444
g2189 and n2442_not n2443_not ; n2445
g2190 and n2444_not n2445_not ; n2446
g2191 and b[24] n266 ; n2447
g2192 and b[22] n284 ; n2448
g2193 and b[23] n261 ; n2449
g2194 and n2448_not n2449_not ; n2450
g2195 and n2447_not n2450 ; n2451
g2196 and n2296_not n2298_not ; n2452
g2197 and b[23]_not b[24]_not ; n2453
g2198 and b[23] b[24] ; n2454
g2199 and n2453_not n2454_not ; n2455
g2200 and n2452_not n2455 ; n2456
g2201 and n2452 n2455_not ; n2457
g2202 and n2456_not n2457_not ; n2458
g2203 and n269 n2458 ; n2459
g2204 and n2451 n2459_not ; n2460
g2205 and a[2] n2460_not ; n2461
g2206 and a[2] n2461_not ; n2462
g2207 and n2460_not n2461_not ; n2463
g2208 and n2462_not n2463_not ; n2464
g2209 and n2446_not n2464_not ; n2465
g2210 and n2446_not n2465_not ; n2466
g2211 and n2464_not n2465_not ; n2467
g2212 and n2466_not n2467_not ; n2468
g2213 and n2307_not n2312_not ; n2469
g2214 and n2468_not n2469_not ; n2470
g2215 and n2468 n2469 ; n2471
g2216 and n2470_not n2471_not ; f[24]
g2217 and n2465_not n2470_not ; n2473
g2218 and b[25] n266 ; n2474
g2219 and b[23] n284 ; n2475
g2220 and b[24] n261 ; n2476
g2221 and n2475_not n2476_not ; n2477
g2222 and n2474_not n2477 ; n2478
g2223 and n2454_not n2456_not ; n2479
g2224 and b[24]_not b[25]_not ; n2480
g2225 and b[24] b[25] ; n2481
g2226 and n2480_not n2481_not ; n2482
g2227 and n2479_not n2482 ; n2483
g2228 and n2479 n2482_not ; n2484
g2229 and n2483_not n2484_not ; n2485
g2230 and n269 n2485 ; n2486
g2231 and n2478 n2486_not ; n2487
g2232 and a[2] n2487_not ; n2488
g2233 and a[2] n2488_not ; n2489
g2234 and n2487_not n2488_not ; n2490
g2235 and n2489_not n2490_not ; n2491
g2236 and n2439_not n2443_not ; n2492
g2237 and b[16] n700 ; n2493
g2238 and b[14] n767 ; n2494
g2239 and b[15] n695 ; n2495
g2240 and n2494_not n2495_not ; n2496
g2241 and n2493_not n2496 ; n2497
g2242 and n703 n1237 ; n2498
g2243 and n2497 n2498_not ; n2499
g2244 and a[11] n2499_not ; n2500
g2245 and a[11] n2500_not ; n2501
g2246 and n2499_not n2500_not ; n2502
g2247 and n2501_not n2502_not ; n2503
g2248 and n2228_not n2387_not ; n2504
g2249 and n2384_not n2504_not ; n2505
g2250 and b[7] n1627 ; n2506
g2251 and b[5] n1763 ; n2507
g2252 and b[6] n1622 ; n2508
g2253 and n2507_not n2508_not ; n2509
g2254 and n2506_not n2509 ; n2510
g2255 and n484 n1630 ; n2511
g2256 and n2510 n2511_not ; n2512
g2257 and a[20] n2512_not ; n2513
g2258 and a[20] n2513_not ; n2514
g2259 and n2512_not n2513_not ; n2515
g2260 and n2514_not n2515_not ; n2516
g2261 and n2210 n2366 ; n2517
g2262 and n2381_not n2517_not ; n2518
g2263 and b[4] n2048 ; n2519
g2264 and b[2] n2198 ; n2520
g2265 and b[3] n2043 ; n2521
g2266 and n2520_not n2521_not ; n2522
g2267 and n2519_not n2522 ; n2523
g2268 and n346 n2051 ; n2524
g2269 and n2523 n2524_not ; n2525
g2270 and a[23] n2525_not ; n2526
g2271 and a[23] n2526_not ; n2527
g2272 and n2525_not n2526_not ; n2528
g2273 and n2527_not n2528_not ; n2529
g2274 and a[26] n2366_not ; n2530
g2275 and a[24]_not a[25] ; n2531
g2276 and a[24] a[25]_not ; n2532
g2277 and n2531_not n2532_not ; n2533
g2278 and n2365 n2533_not ; n2534
g2279 and b[0] n2534 ; n2535
g2280 and a[25]_not a[26] ; n2536
g2281 and a[25] a[26]_not ; n2537
g2282 and n2536_not n2537_not ; n2538
g2283 and n2365_not n2538 ; n2539
g2284 and b[1] n2539 ; n2540
g2285 and n2535_not n2540_not ; n2541
g2286 and n2365_not n2538_not ; n2542
g2287 and n272_not n2542 ; n2543
g2288 and n2541 n2543_not ; n2544
g2289 and a[26] n2544_not ; n2545
g2290 and a[26] n2545_not ; n2546
g2291 and n2544_not n2545_not ; n2547
g2292 and n2546_not n2547_not ; n2548
g2293 and n2530 n2548_not ; n2549
g2294 and n2530_not n2548 ; n2550
g2295 and n2549_not n2550_not ; n2551
g2296 and n2529 n2551 ; n2552
g2297 and n2529_not n2551_not ; n2553
g2298 and n2552_not n2553_not ; n2554
g2299 and n2518_not n2554_not ; n2555
g2300 and n2518 n2554 ; n2556
g2301 and n2555_not n2556_not ; n2557
g2302 and n2516_not n2557 ; n2558
g2303 and n2516 n2557_not ; n2559
g2304 and n2558_not n2559_not ; n2560
g2305 and n2505_not n2560 ; n2561
g2306 and n2505 n2560_not ; n2562
g2307 and n2561_not n2562_not ; n2563
g2308 and b[10] n1302 ; n2564
g2309 and b[8] n1391 ; n2565
g2310 and b[9] n1297 ; n2566
g2311 and n2565_not n2566_not ; n2567
g2312 and n2564_not n2567 ; n2568
g2313 and n738 n1305 ; n2569
g2314 and n2568 n2569_not ; n2570
g2315 and a[17] n2570_not ; n2571
g2316 and a[17] n2571_not ; n2572
g2317 and n2570_not n2571_not ; n2573
g2318 and n2572_not n2573_not ; n2574
g2319 and n2563 n2574_not ; n2575
g2320 and n2563 n2575_not ; n2576
g2321 and n2574_not n2575_not ; n2577
g2322 and n2576_not n2577_not ; n2578
g2323 and n2402_not n2405_not ; n2579
g2324 and n2578 n2579 ; n2580
g2325 and n2578_not n2579_not ; n2581
g2326 and n2580_not n2581_not ; n2582
g2327 and b[13] n951 ; n2583
g2328 and b[11] n1056 ; n2584
g2329 and b[12] n946 ; n2585
g2330 and n2584_not n2585_not ; n2586
g2331 and n2583_not n2586 ; n2587
g2332 and n954 n1008 ; n2588
g2333 and n2587 n2588_not ; n2589
g2334 and a[14] n2589_not ; n2590
g2335 and a[14] n2590_not ; n2591
g2336 and n2589_not n2590_not ; n2592
g2337 and n2591_not n2592_not ; n2593
g2338 and n2582_not n2593 ; n2594
g2339 and n2582 n2593_not ; n2595
g2340 and n2594_not n2595_not ; n2596
g2341 and n2409_not n2411_not ; n2597
g2342 and n2596 n2597_not ; n2598
g2343 and n2596_not n2597 ; n2599
g2344 and n2598_not n2599_not ; n2600
g2345 and n2503_not n2600 ; n2601
g2346 and n2600 n2601_not ; n2602
g2347 and n2503_not n2601_not ; n2603
g2348 and n2602_not n2603_not ; n2604
g2349 and n2414_not n2420_not ; n2605
g2350 and n2604 n2605 ; n2606
g2351 and n2604_not n2605_not ; n2607
g2352 and n2606_not n2607_not ; n2608
g2353 and b[19] n511 ; n2609
g2354 and b[17] n541 ; n2610
g2355 and b[18] n506 ; n2611
g2356 and n2610_not n2611_not ; n2612
g2357 and n2609_not n2612 ; n2613
g2358 and n514 n1708 ; n2614
g2359 and n2613 n2614_not ; n2615
g2360 and a[8] n2615_not ; n2616
g2361 and a[8] n2616_not ; n2617
g2362 and n2615_not n2616_not ; n2618
g2363 and n2617_not n2618_not ; n2619
g2364 and n2608 n2619_not ; n2620
g2365 and n2608 n2620_not ; n2621
g2366 and n2619_not n2620_not ; n2622
g2367 and n2621_not n2622_not ; n2623
g2368 and n2434_not n2436_not ; n2624
g2369 and n2623_not n2624_not ; n2625
g2370 and n2623_not n2625_not ; n2626
g2371 and n2624_not n2625_not ; n2627
g2372 and n2626_not n2627_not ; n2628
g2373 and b[22] n362 ; n2629
g2374 and b[20] n403 ; n2630
g2375 and b[21] n357 ; n2631
g2376 and n2630_not n2631_not ; n2632
g2377 and n2629_not n2632 ; n2633
g2378 and n365 n2145 ; n2634
g2379 and n2633 n2634_not ; n2635
g2380 and a[5] n2635_not ; n2636
g2381 and a[5] n2636_not ; n2637
g2382 and n2635_not n2636_not ; n2638
g2383 and n2637_not n2638_not ; n2639
g2384 and n2628_not n2639 ; n2640
g2385 and n2628 n2639_not ; n2641
g2386 and n2640_not n2641_not ; n2642
g2387 and n2492_not n2642_not ; n2643
g2388 and n2492 n2642 ; n2644
g2389 and n2643_not n2644_not ; n2645
g2390 and n2491_not n2645 ; n2646
g2391 and n2491 n2645_not ; n2647
g2392 and n2646_not n2647_not ; n2648
g2393 and n2473_not n2648 ; n2649
g2394 and n2473 n2648_not ; n2650
g2395 and n2649_not n2650_not ; f[25]
g2396 and n2646_not n2649_not ; n2652
g2397 and n2628_not n2639_not ; n2653
g2398 and n2643_not n2653_not ; n2654
g2399 and n2601_not n2607_not ; n2655
g2400 and n2595_not n2598_not ; n2656
g2401 and b[14] n951 ; n2657
g2402 and b[12] n1056 ; n2658
g2403 and b[13] n946 ; n2659
g2404 and n2658_not n2659_not ; n2660
g2405 and n2657_not n2660 ; n2661
g2406 and n954 n1034 ; n2662
g2407 and n2661 n2662_not ; n2663
g2408 and a[14] n2663_not ; n2664
g2409 and a[14] n2664_not ; n2665
g2410 and n2663_not n2664_not ; n2666
g2411 and n2665_not n2666_not ; n2667
g2412 and n2575_not n2581_not ; n2668
g2413 and b[11] n1302 ; n2669
g2414 and b[9] n1391 ; n2670
g2415 and b[10] n1297 ; n2671
g2416 and n2670_not n2671_not ; n2672
g2417 and n2669_not n2672 ; n2673
g2418 and n818 n1305 ; n2674
g2419 and n2673 n2674_not ; n2675
g2420 and a[17] n2675_not ; n2676
g2421 and a[17] n2676_not ; n2677
g2422 and n2675_not n2676_not ; n2678
g2423 and n2677_not n2678_not ; n2679
g2424 and n2558_not n2561_not ; n2680
g2425 and n2529_not n2551 ; n2681
g2426 and n2555_not n2681_not ; n2682
g2427 and b[2] n2539 ; n2683
g2428 and n2365 n2538_not ; n2684
g2429 and n2533 n2684 ; n2685
g2430 and b[0] n2685 ; n2686
g2431 and b[1] n2534 ; n2687
g2432 and n2686_not n2687_not ; n2688
g2433 and n2683_not n2688 ; n2689
g2434 and n296 n2542 ; n2690
g2435 and n2689 n2690_not ; n2691
g2436 and a[26] n2691_not ; n2692
g2437 and a[26] n2692_not ; n2693
g2438 and n2691_not n2692_not ; n2694
g2439 and n2693_not n2694_not ; n2695
g2440 and n2549_not n2695 ; n2696
g2441 and n2549 n2695_not ; n2697
g2442 and n2696_not n2697_not ; n2698
g2443 and b[5] n2048 ; n2699
g2444 and b[3] n2198 ; n2700
g2445 and b[4] n2043 ; n2701
g2446 and n2700_not n2701_not ; n2702
g2447 and n2699_not n2702 ; n2703
g2448 and n394 n2051 ; n2704
g2449 and n2703 n2704_not ; n2705
g2450 and a[23] n2705_not ; n2706
g2451 and a[23] n2706_not ; n2707
g2452 and n2705_not n2706_not ; n2708
g2453 and n2707_not n2708_not ; n2709
g2454 and n2698 n2709_not ; n2710
g2455 and n2698_not n2709 ; n2711
g2456 and n2682_not n2711_not ; n2712
g2457 and n2710_not n2712 ; n2713
g2458 and n2682_not n2713_not ; n2714
g2459 and n2710_not n2713_not ; n2715
g2460 and n2711_not n2715 ; n2716
g2461 and n2714_not n2716_not ; n2717
g2462 and b[8] n1627 ; n2718
g2463 and b[6] n1763 ; n2719
g2464 and b[7] n1622 ; n2720
g2465 and n2719_not n2720_not ; n2721
g2466 and n2718_not n2721 ; n2722
g2467 and n585 n1630 ; n2723
g2468 and n2722 n2723_not ; n2724
g2469 and a[20] n2724_not ; n2725
g2470 and a[20] n2725_not ; n2726
g2471 and n2724_not n2725_not ; n2727
g2472 and n2726_not n2727_not ; n2728
g2473 and n2717 n2728 ; n2729
g2474 and n2717_not n2728_not ; n2730
g2475 and n2729_not n2730_not ; n2731
g2476 and n2680_not n2731 ; n2732
g2477 and n2680 n2731_not ; n2733
g2478 and n2732_not n2733_not ; n2734
g2479 and n2679 n2734_not ; n2735
g2480 and n2679_not n2734 ; n2736
g2481 and n2735_not n2736_not ; n2737
g2482 and n2668_not n2737 ; n2738
g2483 and n2668 n2737_not ; n2739
g2484 and n2738_not n2739_not ; n2740
g2485 and n2667_not n2740 ; n2741
g2486 and n2740 n2741_not ; n2742
g2487 and n2667_not n2741_not ; n2743
g2488 and n2742_not n2743_not ; n2744
g2489 and n2656_not n2744 ; n2745
g2490 and n2656 n2744_not ; n2746
g2491 and n2745_not n2746_not ; n2747
g2492 and b[17] n700 ; n2748
g2493 and b[15] n767 ; n2749
g2494 and b[16] n695 ; n2750
g2495 and n2749_not n2750_not ; n2751
g2496 and n2748_not n2751 ; n2752
g2497 and n703 n1356 ; n2753
g2498 and n2752 n2753_not ; n2754
g2499 and a[11] n2754_not ; n2755
g2500 and a[11] n2755_not ; n2756
g2501 and n2754_not n2755_not ; n2757
g2502 and n2756_not n2757_not ; n2758
g2503 and n2747_not n2758_not ; n2759
g2504 and n2747 n2758 ; n2760
g2505 and n2759_not n2760_not ; n2761
g2506 and n2655 n2761_not ; n2762
g2507 and n2655_not n2761 ; n2763
g2508 and n2762_not n2763_not ; n2764
g2509 and b[20] n511 ; n2765
g2510 and b[18] n541 ; n2766
g2511 and b[19] n506 ; n2767
g2512 and n2766_not n2767_not ; n2768
g2513 and n2765_not n2768 ; n2769
g2514 and n514 n1846 ; n2770
g2515 and n2769 n2770_not ; n2771
g2516 and a[8] n2771_not ; n2772
g2517 and a[8] n2772_not ; n2773
g2518 and n2771_not n2772_not ; n2774
g2519 and n2773_not n2774_not ; n2775
g2520 and n2764 n2775_not ; n2776
g2521 and n2764 n2776_not ; n2777
g2522 and n2775_not n2776_not ; n2778
g2523 and n2777_not n2778_not ; n2779
g2524 and n2620_not n2625_not ; n2780
g2525 and n2779 n2780 ; n2781
g2526 and n2779_not n2780_not ; n2782
g2527 and n2781_not n2782_not ; n2783
g2528 and b[23] n362 ; n2784
g2529 and b[21] n403 ; n2785
g2530 and b[22] n357 ; n2786
g2531 and n2785_not n2786_not ; n2787
g2532 and n2784_not n2787 ; n2788
g2533 and n365 n2300 ; n2789
g2534 and n2788 n2789_not ; n2790
g2535 and a[5] n2790_not ; n2791
g2536 and a[5] n2791_not ; n2792
g2537 and n2790_not n2791_not ; n2793
g2538 and n2792_not n2793_not ; n2794
g2539 and n2783 n2794_not ; n2795
g2540 and n2783 n2795_not ; n2796
g2541 and n2794_not n2795_not ; n2797
g2542 and n2796_not n2797_not ; n2798
g2543 and n2654_not n2798 ; n2799
g2544 and n2654 n2798_not ; n2800
g2545 and n2799_not n2800_not ; n2801
g2546 and b[26] n266 ; n2802
g2547 and b[24] n284 ; n2803
g2548 and b[25] n261 ; n2804
g2549 and n2803_not n2804_not ; n2805
g2550 and n2802_not n2805 ; n2806
g2551 and n2481_not n2483_not ; n2807
g2552 and b[25]_not b[26]_not ; n2808
g2553 and b[25] b[26] ; n2809
g2554 and n2808_not n2809_not ; n2810
g2555 and n2807_not n2810 ; n2811
g2556 and n2807 n2810_not ; n2812
g2557 and n2811_not n2812_not ; n2813
g2558 and n269 n2813 ; n2814
g2559 and n2806 n2814_not ; n2815
g2560 and a[2] n2815_not ; n2816
g2561 and a[2] n2816_not ; n2817
g2562 and n2815_not n2816_not ; n2818
g2563 and n2817_not n2818_not ; n2819
g2564 and n2801_not n2819_not ; n2820
g2565 and n2801 n2819 ; n2821
g2566 and n2820_not n2821_not ; n2822
g2567 and n2652_not n2822 ; n2823
g2568 and n2652 n2822_not ; n2824
g2569 and n2823_not n2824_not ; f[26]
g2570 and n2820_not n2823_not ; n2826
g2571 and b[24] n362 ; n2827
g2572 and b[22] n403 ; n2828
g2573 and b[23] n357 ; n2829
g2574 and n2828_not n2829_not ; n2830
g2575 and n2827_not n2830 ; n2831
g2576 and n365 n2458 ; n2832
g2577 and n2831 n2832_not ; n2833
g2578 and a[5] n2833_not ; n2834
g2579 and a[5] n2834_not ; n2835
g2580 and n2833_not n2834_not ; n2836
g2581 and n2835_not n2836_not ; n2837
g2582 and b[15] n951 ; n2838
g2583 and b[13] n1056 ; n2839
g2584 and b[14] n946 ; n2840
g2585 and n2839_not n2840_not ; n2841
g2586 and n2838_not n2841 ; n2842
g2587 and n954 n1131 ; n2843
g2588 and n2842 n2843_not ; n2844
g2589 and a[14] n2844_not ; n2845
g2590 and a[14] n2845_not ; n2846
g2591 and n2844_not n2845_not ; n2847
g2592 and n2846_not n2847_not ; n2848
g2593 and n2736_not n2738_not ; n2849
g2594 and b[12] n1302 ; n2850
g2595 and b[10] n1391 ; n2851
g2596 and b[11] n1297 ; n2852
g2597 and n2851_not n2852_not ; n2853
g2598 and n2850_not n2853 ; n2854
g2599 and n842 n1305 ; n2855
g2600 and n2854 n2855_not ; n2856
g2601 and a[17] n2856_not ; n2857
g2602 and a[17] n2857_not ; n2858
g2603 and n2856_not n2857_not ; n2859
g2604 and n2858_not n2859_not ; n2860
g2605 and n2730_not n2732_not ; n2861
g2606 and b[6] n2048 ; n2862
g2607 and b[4] n2198 ; n2863
g2608 and b[5] n2043 ; n2864
g2609 and n2863_not n2864_not ; n2865
g2610 and n2862_not n2865 ; n2866
g2611 and n459 n2051 ; n2867
g2612 and n2866 n2867_not ; n2868
g2613 and a[23] n2868_not ; n2869
g2614 and a[23] n2869_not ; n2870
g2615 and n2868_not n2869_not ; n2871
g2616 and n2870_not n2871_not ; n2872
g2617 and a[26] a[27]_not ; n2873
g2618 and a[26]_not a[27] ; n2874
g2619 and n2873_not n2874_not ; n2875
g2620 and b[0] n2875_not ; n2876
g2621 and n2697_not n2876 ; n2877
g2622 and n2697 n2876_not ; n2878
g2623 and n2877_not n2878_not ; n2879
g2624 and b[3] n2539 ; n2880
g2625 and b[1] n2685 ; n2881
g2626 and b[2] n2534 ; n2882
g2627 and n2881_not n2882_not ; n2883
g2628 and n2880_not n2883 ; n2884
g2629 and n318 n2542 ; n2885
g2630 and n2884 n2885_not ; n2886
g2631 and a[26] n2886_not ; n2887
g2632 and a[26] n2887_not ; n2888
g2633 and n2886_not n2887_not ; n2889
g2634 and n2888_not n2889_not ; n2890
g2635 and n2879_not n2890_not ; n2891
g2636 and n2879 n2890 ; n2892
g2637 and n2891_not n2892_not ; n2893
g2638 and n2872_not n2893 ; n2894
g2639 and n2893 n2894_not ; n2895
g2640 and n2872_not n2894_not ; n2896
g2641 and n2895_not n2896_not ; n2897
g2642 and n2715_not n2897 ; n2898
g2643 and n2715 n2897_not ; n2899
g2644 and n2898_not n2899_not ; n2900
g2645 and b[9] n1627 ; n2901
g2646 and b[7] n1763 ; n2902
g2647 and b[8] n1622 ; n2903
g2648 and n2902_not n2903_not ; n2904
g2649 and n2901_not n2904 ; n2905
g2650 and n651 n1630 ; n2906
g2651 and n2905 n2906_not ; n2907
g2652 and a[20] n2907_not ; n2908
g2653 and a[20] n2908_not ; n2909
g2654 and n2907_not n2908_not ; n2910
g2655 and n2909_not n2910_not ; n2911
g2656 and n2900_not n2911_not ; n2912
g2657 and n2900 n2911 ; n2913
g2658 and n2912_not n2913_not ; n2914
g2659 and n2861_not n2914 ; n2915
g2660 and n2861 n2914_not ; n2916
g2661 and n2915_not n2916_not ; n2917
g2662 and n2860 n2917_not ; n2918
g2663 and n2860_not n2917 ; n2919
g2664 and n2918_not n2919_not ; n2920
g2665 and n2849_not n2920 ; n2921
g2666 and n2849 n2920_not ; n2922
g2667 and n2921_not n2922_not ; n2923
g2668 and n2848_not n2923 ; n2924
g2669 and n2923 n2924_not ; n2925
g2670 and n2848_not n2924_not ; n2926
g2671 and n2925_not n2926_not ; n2927
g2672 and n2656_not n2744_not ; n2928
g2673 and n2741_not n2928_not ; n2929
g2674 and n2927 n2929 ; n2930
g2675 and n2927_not n2929_not ; n2931
g2676 and n2930_not n2931_not ; n2932
g2677 and b[18] n700 ; n2933
g2678 and b[16] n767 ; n2934
g2679 and b[17] n695 ; n2935
g2680 and n2934_not n2935_not ; n2936
g2681 and n2933_not n2936 ; n2937
g2682 and n703 n1566 ; n2938
g2683 and n2937 n2938_not ; n2939
g2684 and a[11] n2939_not ; n2940
g2685 and a[11] n2940_not ; n2941
g2686 and n2939_not n2940_not ; n2942
g2687 and n2941_not n2942_not ; n2943
g2688 and n2932 n2943_not ; n2944
g2689 and n2932 n2944_not ; n2945
g2690 and n2943_not n2944_not ; n2946
g2691 and n2945_not n2946_not ; n2947
g2692 and n2759_not n2763_not ; n2948
g2693 and n2947 n2948 ; n2949
g2694 and n2947_not n2948_not ; n2950
g2695 and n2949_not n2950_not ; n2951
g2696 and b[21] n511 ; n2952
g2697 and b[19] n541 ; n2953
g2698 and b[20] n506 ; n2954
g2699 and n2953_not n2954_not ; n2955
g2700 and n2952_not n2955 ; n2956
g2701 and n514 n1984 ; n2957
g2702 and n2956 n2957_not ; n2958
g2703 and a[8] n2958_not ; n2959
g2704 and a[8] n2959_not ; n2960
g2705 and n2958_not n2959_not ; n2961
g2706 and n2960_not n2961_not ; n2962
g2707 and n2951_not n2962 ; n2963
g2708 and n2951 n2962_not ; n2964
g2709 and n2963_not n2964_not ; n2965
g2710 and n2776_not n2782_not ; n2966
g2711 and n2965 n2966_not ; n2967
g2712 and n2965_not n2966 ; n2968
g2713 and n2967_not n2968_not ; n2969
g2714 and n2837_not n2969 ; n2970
g2715 and n2969 n2970_not ; n2971
g2716 and n2837_not n2970_not ; n2972
g2717 and n2971_not n2972_not ; n2973
g2718 and n2654_not n2798_not ; n2974
g2719 and n2795_not n2974_not ; n2975
g2720 and n2973 n2975 ; n2976
g2721 and n2973_not n2975_not ; n2977
g2722 and n2976_not n2977_not ; n2978
g2723 and b[27] n266 ; n2979
g2724 and b[25] n284 ; n2980
g2725 and b[26] n261 ; n2981
g2726 and n2980_not n2981_not ; n2982
g2727 and n2979_not n2982 ; n2983
g2728 and n2809_not n2811_not ; n2984
g2729 and b[26]_not b[27]_not ; n2985
g2730 and b[26] b[27] ; n2986
g2731 and n2985_not n2986_not ; n2987
g2732 and n2984_not n2987 ; n2988
g2733 and n2984 n2987_not ; n2989
g2734 and n2988_not n2989_not ; n2990
g2735 and n269 n2990 ; n2991
g2736 and n2983 n2991_not ; n2992
g2737 and a[2] n2992_not ; n2993
g2738 and a[2] n2993_not ; n2994
g2739 and n2992_not n2993_not ; n2995
g2740 and n2994_not n2995_not ; n2996
g2741 and n2978_not n2996 ; n2997
g2742 and n2978 n2996_not ; n2998
g2743 and n2997_not n2998_not ; n2999
g2744 and n2826_not n2999 ; n3000
g2745 and n2826 n2999_not ; n3001
g2746 and n3000_not n3001_not ; f[27]
g2747 and n2998_not n3000_not ; n3003
g2748 and b[25] n362 ; n3004
g2749 and b[23] n403 ; n3005
g2750 and b[24] n357 ; n3006
g2751 and n3005_not n3006_not ; n3007
g2752 and n3004_not n3007 ; n3008
g2753 and n365 n2485 ; n3009
g2754 and n3008 n3009_not ; n3010
g2755 and a[5] n3010_not ; n3011
g2756 and a[5] n3011_not ; n3012
g2757 and n3010_not n3011_not ; n3013
g2758 and n3012_not n3013_not ; n3014
g2759 and n2715_not n2897_not ; n3015
g2760 and n2894_not n3015_not ; n3016
g2761 and b[7] n2048 ; n3017
g2762 and b[5] n2198 ; n3018
g2763 and b[6] n2043 ; n3019
g2764 and n3018_not n3019_not ; n3020
g2765 and n3017_not n3020 ; n3021
g2766 and n484 n2051 ; n3022
g2767 and n3021 n3022_not ; n3023
g2768 and a[23] n3023_not ; n3024
g2769 and a[23] n3024_not ; n3025
g2770 and n3023_not n3024_not ; n3026
g2771 and n3025_not n3026_not ; n3027
g2772 and n2697 n2876 ; n3028
g2773 and n2891_not n3028_not ; n3029
g2774 and b[4] n2539 ; n3030
g2775 and b[2] n2685 ; n3031
g2776 and b[3] n2534 ; n3032
g2777 and n3031_not n3032_not ; n3033
g2778 and n3030_not n3033 ; n3034
g2779 and n346 n2542 ; n3035
g2780 and n3034 n3035_not ; n3036
g2781 and a[26] n3036_not ; n3037
g2782 and a[26] n3037_not ; n3038
g2783 and n3036_not n3037_not ; n3039
g2784 and n3038_not n3039_not ; n3040
g2785 and a[29] n2876_not ; n3041
g2786 and a[27]_not a[28] ; n3042
g2787 and a[27] a[28]_not ; n3043
g2788 and n3042_not n3043_not ; n3044
g2789 and n2875 n3044_not ; n3045
g2790 and b[0] n3045 ; n3046
g2791 and a[28]_not a[29] ; n3047
g2792 and a[28] a[29]_not ; n3048
g2793 and n3047_not n3048_not ; n3049
g2794 and n2875_not n3049 ; n3050
g2795 and b[1] n3050 ; n3051
g2796 and n3046_not n3051_not ; n3052
g2797 and n2875_not n3049_not ; n3053
g2798 and n272_not n3053 ; n3054
g2799 and n3052 n3054_not ; n3055
g2800 and a[29] n3055_not ; n3056
g2801 and a[29] n3056_not ; n3057
g2802 and n3055_not n3056_not ; n3058
g2803 and n3057_not n3058_not ; n3059
g2804 and n3041 n3059_not ; n3060
g2805 and n3041_not n3059 ; n3061
g2806 and n3060_not n3061_not ; n3062
g2807 and n3040 n3062 ; n3063
g2808 and n3040_not n3062_not ; n3064
g2809 and n3063_not n3064_not ; n3065
g2810 and n3029_not n3065_not ; n3066
g2811 and n3029 n3065 ; n3067
g2812 and n3066_not n3067_not ; n3068
g2813 and n3027_not n3068 ; n3069
g2814 and n3027 n3068_not ; n3070
g2815 and n3069_not n3070_not ; n3071
g2816 and n3016_not n3071 ; n3072
g2817 and n3016 n3071_not ; n3073
g2818 and n3072_not n3073_not ; n3074
g2819 and b[10] n1627 ; n3075
g2820 and b[8] n1763 ; n3076
g2821 and b[9] n1622 ; n3077
g2822 and n3076_not n3077_not ; n3078
g2823 and n3075_not n3078 ; n3079
g2824 and n738 n1630 ; n3080
g2825 and n3079 n3080_not ; n3081
g2826 and a[20] n3081_not ; n3082
g2827 and a[20] n3082_not ; n3083
g2828 and n3081_not n3082_not ; n3084
g2829 and n3083_not n3084_not ; n3085
g2830 and n3074 n3085_not ; n3086
g2831 and n3074 n3086_not ; n3087
g2832 and n3085_not n3086_not ; n3088
g2833 and n3087_not n3088_not ; n3089
g2834 and n2912_not n2915_not ; n3090
g2835 and n3089 n3090 ; n3091
g2836 and n3089_not n3090_not ; n3092
g2837 and n3091_not n3092_not ; n3093
g2838 and b[13] n1302 ; n3094
g2839 and b[11] n1391 ; n3095
g2840 and b[12] n1297 ; n3096
g2841 and n3095_not n3096_not ; n3097
g2842 and n3094_not n3097 ; n3098
g2843 and n1008 n1305 ; n3099
g2844 and n3098 n3099_not ; n3100
g2845 and a[17] n3100_not ; n3101
g2846 and a[17] n3101_not ; n3102
g2847 and n3100_not n3101_not ; n3103
g2848 and n3102_not n3103_not ; n3104
g2849 and n3093 n3104_not ; n3105
g2850 and n3093 n3105_not ; n3106
g2851 and n3104_not n3105_not ; n3107
g2852 and n3106_not n3107_not ; n3108
g2853 and n2919_not n2921_not ; n3109
g2854 and n3108_not n3109_not ; n3110
g2855 and n3108_not n3110_not ; n3111
g2856 and n3109_not n3110_not ; n3112
g2857 and n3111_not n3112_not ; n3113
g2858 and b[16] n951 ; n3114
g2859 and b[14] n1056 ; n3115
g2860 and b[15] n946 ; n3116
g2861 and n3115_not n3116_not ; n3117
g2862 and n3114_not n3117 ; n3118
g2863 and n954 n1237 ; n3119
g2864 and n3118 n3119_not ; n3120
g2865 and a[14] n3120_not ; n3121
g2866 and a[14] n3121_not ; n3122
g2867 and n3120_not n3121_not ; n3123
g2868 and n3122_not n3123_not ; n3124
g2869 and n3113_not n3124_not ; n3125
g2870 and n3113_not n3125_not ; n3126
g2871 and n3124_not n3125_not ; n3127
g2872 and n3126_not n3127_not ; n3128
g2873 and n2924_not n2931_not ; n3129
g2874 and n3128 n3129 ; n3130
g2875 and n3128_not n3129_not ; n3131
g2876 and n3130_not n3131_not ; n3132
g2877 and b[19] n700 ; n3133
g2878 and b[17] n767 ; n3134
g2879 and b[18] n695 ; n3135
g2880 and n3134_not n3135_not ; n3136
g2881 and n3133_not n3136 ; n3137
g2882 and n703 n1708 ; n3138
g2883 and n3137 n3138_not ; n3139
g2884 and a[11] n3139_not ; n3140
g2885 and a[11] n3140_not ; n3141
g2886 and n3139_not n3140_not ; n3142
g2887 and n3141_not n3142_not ; n3143
g2888 and n3132 n3143_not ; n3144
g2889 and n3132 n3144_not ; n3145
g2890 and n3143_not n3144_not ; n3146
g2891 and n3145_not n3146_not ; n3147
g2892 and n2944_not n2950_not ; n3148
g2893 and n3147 n3148 ; n3149
g2894 and n3147_not n3148_not ; n3150
g2895 and n3149_not n3150_not ; n3151
g2896 and b[22] n511 ; n3152
g2897 and b[20] n541 ; n3153
g2898 and b[21] n506 ; n3154
g2899 and n3153_not n3154_not ; n3155
g2900 and n3152_not n3155 ; n3156
g2901 and n514 n2145 ; n3157
g2902 and n3156 n3157_not ; n3158
g2903 and a[8] n3158_not ; n3159
g2904 and a[8] n3159_not ; n3160
g2905 and n3158_not n3159_not ; n3161
g2906 and n3160_not n3161_not ; n3162
g2907 and n3151_not n3162 ; n3163
g2908 and n3151 n3162_not ; n3164
g2909 and n3163_not n3164_not ; n3165
g2910 and n2964_not n2967_not ; n3166
g2911 and n3165 n3166_not ; n3167
g2912 and n3165_not n3166 ; n3168
g2913 and n3167_not n3168_not ; n3169
g2914 and n3014_not n3169 ; n3170
g2915 and n3169 n3170_not ; n3171
g2916 and n3014_not n3170_not ; n3172
g2917 and n3171_not n3172_not ; n3173
g2918 and n2970_not n2977_not ; n3174
g2919 and n3173 n3174 ; n3175
g2920 and n3173_not n3174_not ; n3176
g2921 and n3175_not n3176_not ; n3177
g2922 and b[28] n266 ; n3178
g2923 and b[26] n284 ; n3179
g2924 and b[27] n261 ; n3180
g2925 and n3179_not n3180_not ; n3181
g2926 and n3178_not n3181 ; n3182
g2927 and n2986_not n2988_not ; n3183
g2928 and b[27]_not b[28]_not ; n3184
g2929 and b[27] b[28] ; n3185
g2930 and n3184_not n3185_not ; n3186
g2931 and n3183_not n3186 ; n3187
g2932 and n3183 n3186_not ; n3188
g2933 and n3187_not n3188_not ; n3189
g2934 and n269 n3189 ; n3190
g2935 and n3182 n3190_not ; n3191
g2936 and a[2] n3191_not ; n3192
g2937 and a[2] n3192_not ; n3193
g2938 and n3191_not n3192_not ; n3194
g2939 and n3193_not n3194_not ; n3195
g2940 and n3177_not n3195 ; n3196
g2941 and n3177 n3195_not ; n3197
g2942 and n3196_not n3197_not ; n3198
g2943 and n3003_not n3198 ; n3199
g2944 and n3003 n3198_not ; n3200
g2945 and n3199_not n3200_not ; f[28]
g2946 and n3170_not n3176_not ; n3202
g2947 and b[26] n362 ; n3203
g2948 and b[24] n403 ; n3204
g2949 and b[25] n357 ; n3205
g2950 and n3204_not n3205_not ; n3206
g2951 and n3203_not n3206 ; n3207
g2952 and n365 n2813 ; n3208
g2953 and n3207 n3208_not ; n3209
g2954 and a[5] n3209_not ; n3210
g2955 and a[5] n3210_not ; n3211
g2956 and n3209_not n3210_not ; n3212
g2957 and n3211_not n3212_not ; n3213
g2958 and n3144_not n3150_not ; n3214
g2959 and b[14] n1302 ; n3215
g2960 and b[12] n1391 ; n3216
g2961 and b[13] n1297 ; n3217
g2962 and n3216_not n3217_not ; n3218
g2963 and n3215_not n3218 ; n3219
g2964 and n1034 n1305 ; n3220
g2965 and n3219 n3220_not ; n3221
g2966 and a[17] n3221_not ; n3222
g2967 and a[17] n3222_not ; n3223
g2968 and n3221_not n3222_not ; n3224
g2969 and n3223_not n3224_not ; n3225
g2970 and n3086_not n3092_not ; n3226
g2971 and b[11] n1627 ; n3227
g2972 and b[9] n1763 ; n3228
g2973 and b[10] n1622 ; n3229
g2974 and n3228_not n3229_not ; n3230
g2975 and n3227_not n3230 ; n3231
g2976 and n818 n1630 ; n3232
g2977 and n3231 n3232_not ; n3233
g2978 and a[20] n3233_not ; n3234
g2979 and a[20] n3234_not ; n3235
g2980 and n3233_not n3234_not ; n3236
g2981 and n3235_not n3236_not ; n3237
g2982 and n3069_not n3072_not ; n3238
g2983 and n3040_not n3062 ; n3239
g2984 and n3066_not n3239_not ; n3240
g2985 and b[2] n3050 ; n3241
g2986 and n2875 n3049_not ; n3242
g2987 and n3044 n3242 ; n3243
g2988 and b[0] n3243 ; n3244
g2989 and b[1] n3045 ; n3245
g2990 and n3244_not n3245_not ; n3246
g2991 and n3241_not n3246 ; n3247
g2992 and n296 n3053 ; n3248
g2993 and n3247 n3248_not ; n3249
g2994 and a[29] n3249_not ; n3250
g2995 and a[29] n3250_not ; n3251
g2996 and n3249_not n3250_not ; n3252
g2997 and n3251_not n3252_not ; n3253
g2998 and n3060_not n3253 ; n3254
g2999 and n3060 n3253_not ; n3255
g3000 and n3254_not n3255_not ; n3256
g3001 and b[5] n2539 ; n3257
g3002 and b[3] n2685 ; n3258
g3003 and b[4] n2534 ; n3259
g3004 and n3258_not n3259_not ; n3260
g3005 and n3257_not n3260 ; n3261
g3006 and n394 n2542 ; n3262
g3007 and n3261 n3262_not ; n3263
g3008 and a[26] n3263_not ; n3264
g3009 and a[26] n3264_not ; n3265
g3010 and n3263_not n3264_not ; n3266
g3011 and n3265_not n3266_not ; n3267
g3012 and n3256 n3267_not ; n3268
g3013 and n3256_not n3267 ; n3269
g3014 and n3240_not n3269_not ; n3270
g3015 and n3268_not n3270 ; n3271
g3016 and n3240_not n3271_not ; n3272
g3017 and n3268_not n3271_not ; n3273
g3018 and n3269_not n3273 ; n3274
g3019 and n3272_not n3274_not ; n3275
g3020 and b[8] n2048 ; n3276
g3021 and b[6] n2198 ; n3277
g3022 and b[7] n2043 ; n3278
g3023 and n3277_not n3278_not ; n3279
g3024 and n3276_not n3279 ; n3280
g3025 and n585 n2051 ; n3281
g3026 and n3280 n3281_not ; n3282
g3027 and a[23] n3282_not ; n3283
g3028 and a[23] n3283_not ; n3284
g3029 and n3282_not n3283_not ; n3285
g3030 and n3284_not n3285_not ; n3286
g3031 and n3275 n3286 ; n3287
g3032 and n3275_not n3286_not ; n3288
g3033 and n3287_not n3288_not ; n3289
g3034 and n3238_not n3289 ; n3290
g3035 and n3238 n3289_not ; n3291
g3036 and n3290_not n3291_not ; n3292
g3037 and n3237 n3292_not ; n3293
g3038 and n3237_not n3292 ; n3294
g3039 and n3293_not n3294_not ; n3295
g3040 and n3226_not n3295 ; n3296
g3041 and n3226 n3295_not ; n3297
g3042 and n3296_not n3297_not ; n3298
g3043 and n3225_not n3298 ; n3299
g3044 and n3298 n3299_not ; n3300
g3045 and n3225_not n3299_not ; n3301
g3046 and n3300_not n3301_not ; n3302
g3047 and n3105_not n3110_not ; n3303
g3048 and n3302 n3303 ; n3304
g3049 and n3302_not n3303_not ; n3305
g3050 and n3304_not n3305_not ; n3306
g3051 and b[17] n951 ; n3307
g3052 and b[15] n1056 ; n3308
g3053 and b[16] n946 ; n3309
g3054 and n3308_not n3309_not ; n3310
g3055 and n3307_not n3310 ; n3311
g3056 and n954 n1356 ; n3312
g3057 and n3311 n3312_not ; n3313
g3058 and a[14] n3313_not ; n3314
g3059 and a[14] n3314_not ; n3315
g3060 and n3313_not n3314_not ; n3316
g3061 and n3315_not n3316_not ; n3317
g3062 and n3306 n3317_not ; n3318
g3063 and n3306 n3318_not ; n3319
g3064 and n3317_not n3318_not ; n3320
g3065 and n3319_not n3320_not ; n3321
g3066 and n3125_not n3131_not ; n3322
g3067 and n3321 n3322 ; n3323
g3068 and n3321_not n3322_not ; n3324
g3069 and n3323_not n3324_not ; n3325
g3070 and b[20] n700 ; n3326
g3071 and b[18] n767 ; n3327
g3072 and b[19] n695 ; n3328
g3073 and n3327_not n3328_not ; n3329
g3074 and n3326_not n3329 ; n3330
g3075 and n703 n1846 ; n3331
g3076 and n3330 n3331_not ; n3332
g3077 and a[11] n3332_not ; n3333
g3078 and a[11] n3333_not ; n3334
g3079 and n3332_not n3333_not ; n3335
g3080 and n3334_not n3335_not ; n3336
g3081 and n3325 n3336_not ; n3337
g3082 and n3325_not n3336 ; n3338
g3083 and n3214_not n3338_not ; n3339
g3084 and n3337_not n3339 ; n3340
g3085 and n3214_not n3340_not ; n3341
g3086 and n3337_not n3340_not ; n3342
g3087 and n3338_not n3342 ; n3343
g3088 and n3341_not n3343_not ; n3344
g3089 and b[23] n511 ; n3345
g3090 and b[21] n541 ; n3346
g3091 and b[22] n506 ; n3347
g3092 and n3346_not n3347_not ; n3348
g3093 and n3345_not n3348 ; n3349
g3094 and n514 n2300 ; n3350
g3095 and n3349 n3350_not ; n3351
g3096 and a[8] n3351_not ; n3352
g3097 and a[8] n3352_not ; n3353
g3098 and n3351_not n3352_not ; n3354
g3099 and n3353_not n3354_not ; n3355
g3100 and n3344_not n3355_not ; n3356
g3101 and n3344_not n3356_not ; n3357
g3102 and n3355_not n3356_not ; n3358
g3103 and n3357_not n3358_not ; n3359
g3104 and n3164_not n3167_not ; n3360
g3105 and n3359_not n3360_not ; n3361
g3106 and n3359 n3360 ; n3362
g3107 and n3361_not n3362_not ; n3363
g3108 and n3213_not n3363 ; n3364
g3109 and n3213_not n3364_not ; n3365
g3110 and n3363 n3364_not ; n3366
g3111 and n3365_not n3366_not ; n3367
g3112 and n3202_not n3367_not ; n3368
g3113 and n3202_not n3368_not ; n3369
g3114 and n3367_not n3368_not ; n3370
g3115 and n3369_not n3370_not ; n3371
g3116 and b[29] n266 ; n3372
g3117 and b[27] n284 ; n3373
g3118 and b[28] n261 ; n3374
g3119 and n3373_not n3374_not ; n3375
g3120 and n3372_not n3375 ; n3376
g3121 and n3185_not n3187_not ; n3377
g3122 and b[28]_not b[29]_not ; n3378
g3123 and b[28] b[29] ; n3379
g3124 and n3378_not n3379_not ; n3380
g3125 and n3377_not n3380 ; n3381
g3126 and n3377 n3380_not ; n3382
g3127 and n3381_not n3382_not ; n3383
g3128 and n269 n3383 ; n3384
g3129 and n3376 n3384_not ; n3385
g3130 and a[2] n3385_not ; n3386
g3131 and a[2] n3386_not ; n3387
g3132 and n3385_not n3386_not ; n3388
g3133 and n3387_not n3388_not ; n3389
g3134 and n3371_not n3389_not ; n3390
g3135 and n3371_not n3390_not ; n3391
g3136 and n3389_not n3390_not ; n3392
g3137 and n3391_not n3392_not ; n3393
g3138 and n3197_not n3199_not ; n3394
g3139 and n3393_not n3394_not ; n3395
g3140 and n3393 n3394 ; n3396
g3141 and n3395_not n3396_not ; f[29]
g3142 and n3356_not n3361_not ; n3398
g3143 and b[15] n1302 ; n3399
g3144 and b[13] n1391 ; n3400
g3145 and b[14] n1297 ; n3401
g3146 and n3400_not n3401_not ; n3402
g3147 and n3399_not n3402 ; n3403
g3148 and n1131 n1305 ; n3404
g3149 and n3403 n3404_not ; n3405
g3150 and a[17] n3405_not ; n3406
g3151 and a[17] n3406_not ; n3407
g3152 and n3405_not n3406_not ; n3408
g3153 and n3407_not n3408_not ; n3409
g3154 and n3294_not n3296_not ; n3410
g3155 and b[12] n1627 ; n3411
g3156 and b[10] n1763 ; n3412
g3157 and b[11] n1622 ; n3413
g3158 and n3412_not n3413_not ; n3414
g3159 and n3411_not n3414 ; n3415
g3160 and n842 n1630 ; n3416
g3161 and n3415 n3416_not ; n3417
g3162 and a[20] n3417_not ; n3418
g3163 and a[20] n3418_not ; n3419
g3164 and n3417_not n3418_not ; n3420
g3165 and n3419_not n3420_not ; n3421
g3166 and n3288_not n3290_not ; n3422
g3167 and b[6] n2539 ; n3423
g3168 and b[4] n2685 ; n3424
g3169 and b[5] n2534 ; n3425
g3170 and n3424_not n3425_not ; n3426
g3171 and n3423_not n3426 ; n3427
g3172 and n459 n2542 ; n3428
g3173 and n3427 n3428_not ; n3429
g3174 and a[26] n3429_not ; n3430
g3175 and a[26] n3430_not ; n3431
g3176 and n3429_not n3430_not ; n3432
g3177 and n3431_not n3432_not ; n3433
g3178 and a[29] a[30]_not ; n3434
g3179 and a[29]_not a[30] ; n3435
g3180 and n3434_not n3435_not ; n3436
g3181 and b[0] n3436_not ; n3437
g3182 and n3255_not n3437 ; n3438
g3183 and n3255 n3437_not ; n3439
g3184 and n3438_not n3439_not ; n3440
g3185 and b[3] n3050 ; n3441
g3186 and b[1] n3243 ; n3442
g3187 and b[2] n3045 ; n3443
g3188 and n3442_not n3443_not ; n3444
g3189 and n3441_not n3444 ; n3445
g3190 and n318 n3053 ; n3446
g3191 and n3445 n3446_not ; n3447
g3192 and a[29] n3447_not ; n3448
g3193 and a[29] n3448_not ; n3449
g3194 and n3447_not n3448_not ; n3450
g3195 and n3449_not n3450_not ; n3451
g3196 and n3440_not n3451_not ; n3452
g3197 and n3440 n3451 ; n3453
g3198 and n3452_not n3453_not ; n3454
g3199 and n3433_not n3454 ; n3455
g3200 and n3454 n3455_not ; n3456
g3201 and n3433_not n3455_not ; n3457
g3202 and n3456_not n3457_not ; n3458
g3203 and n3273_not n3458 ; n3459
g3204 and n3273 n3458_not ; n3460
g3205 and n3459_not n3460_not ; n3461
g3206 and b[9] n2048 ; n3462
g3207 and b[7] n2198 ; n3463
g3208 and b[8] n2043 ; n3464
g3209 and n3463_not n3464_not ; n3465
g3210 and n3462_not n3465 ; n3466
g3211 and n651 n2051 ; n3467
g3212 and n3466 n3467_not ; n3468
g3213 and a[23] n3468_not ; n3469
g3214 and a[23] n3469_not ; n3470
g3215 and n3468_not n3469_not ; n3471
g3216 and n3470_not n3471_not ; n3472
g3217 and n3461_not n3472_not ; n3473
g3218 and n3461 n3472 ; n3474
g3219 and n3473_not n3474_not ; n3475
g3220 and n3422_not n3475 ; n3476
g3221 and n3422 n3475_not ; n3477
g3222 and n3476_not n3477_not ; n3478
g3223 and n3421 n3478_not ; n3479
g3224 and n3421_not n3478 ; n3480
g3225 and n3479_not n3480_not ; n3481
g3226 and n3410_not n3481 ; n3482
g3227 and n3410 n3481_not ; n3483
g3228 and n3482_not n3483_not ; n3484
g3229 and n3409_not n3484 ; n3485
g3230 and n3484 n3485_not ; n3486
g3231 and n3409_not n3485_not ; n3487
g3232 and n3486_not n3487_not ; n3488
g3233 and n3299_not n3305_not ; n3489
g3234 and n3488 n3489 ; n3490
g3235 and n3488_not n3489_not ; n3491
g3236 and n3490_not n3491_not ; n3492
g3237 and b[18] n951 ; n3493
g3238 and b[16] n1056 ; n3494
g3239 and b[17] n946 ; n3495
g3240 and n3494_not n3495_not ; n3496
g3241 and n3493_not n3496 ; n3497
g3242 and n954 n1566 ; n3498
g3243 and n3497 n3498_not ; n3499
g3244 and a[14] n3499_not ; n3500
g3245 and a[14] n3500_not ; n3501
g3246 and n3499_not n3500_not ; n3502
g3247 and n3501_not n3502_not ; n3503
g3248 and n3492 n3503_not ; n3504
g3249 and n3492 n3504_not ; n3505
g3250 and n3503_not n3504_not ; n3506
g3251 and n3505_not n3506_not ; n3507
g3252 and n3318_not n3324_not ; n3508
g3253 and n3507 n3508 ; n3509
g3254 and n3507_not n3508_not ; n3510
g3255 and n3509_not n3510_not ; n3511
g3256 and b[21] n700 ; n3512
g3257 and b[19] n767 ; n3513
g3258 and b[20] n695 ; n3514
g3259 and n3513_not n3514_not ; n3515
g3260 and n3512_not n3515 ; n3516
g3261 and n703 n1984 ; n3517
g3262 and n3516 n3517_not ; n3518
g3263 and a[11] n3518_not ; n3519
g3264 and a[11] n3519_not ; n3520
g3265 and n3518_not n3519_not ; n3521
g3266 and n3520_not n3521_not ; n3522
g3267 and n3511 n3522_not ; n3523
g3268 and n3511 n3523_not ; n3524
g3269 and n3522_not n3523_not ; n3525
g3270 and n3524_not n3525_not ; n3526
g3271 and n3342_not n3526 ; n3527
g3272 and n3342 n3526_not ; n3528
g3273 and n3527_not n3528_not ; n3529
g3274 and b[24] n511 ; n3530
g3275 and b[22] n541 ; n3531
g3276 and b[23] n506 ; n3532
g3277 and n3531_not n3532_not ; n3533
g3278 and n3530_not n3533 ; n3534
g3279 and n514 n2458 ; n3535
g3280 and n3534 n3535_not ; n3536
g3281 and a[8] n3536_not ; n3537
g3282 and a[8] n3537_not ; n3538
g3283 and n3536_not n3537_not ; n3539
g3284 and n3538_not n3539_not ; n3540
g3285 and n3529_not n3540_not ; n3541
g3286 and n3529 n3540 ; n3542
g3287 and n3541_not n3542_not ; n3543
g3288 and n3398 n3543_not ; n3544
g3289 and n3398_not n3543 ; n3545
g3290 and n3544_not n3545_not ; n3546
g3291 and b[27] n362 ; n3547
g3292 and b[25] n403 ; n3548
g3293 and b[26] n357 ; n3549
g3294 and n3548_not n3549_not ; n3550
g3295 and n3547_not n3550 ; n3551
g3296 and n365 n2990 ; n3552
g3297 and n3551 n3552_not ; n3553
g3298 and a[5] n3553_not ; n3554
g3299 and a[5] n3554_not ; n3555
g3300 and n3553_not n3554_not ; n3556
g3301 and n3555_not n3556_not ; n3557
g3302 and n3546 n3557_not ; n3558
g3303 and n3546 n3558_not ; n3559
g3304 and n3557_not n3558_not ; n3560
g3305 and n3559_not n3560_not ; n3561
g3306 and n3364_not n3368_not ; n3562
g3307 and n3561 n3562 ; n3563
g3308 and n3561_not n3562_not ; n3564
g3309 and n3563_not n3564_not ; n3565
g3310 and b[30] n266 ; n3566
g3311 and b[28] n284 ; n3567
g3312 and b[29] n261 ; n3568
g3313 and n3567_not n3568_not ; n3569
g3314 and n3566_not n3569 ; n3570
g3315 and n3379_not n3381_not ; n3571
g3316 and b[29]_not b[30]_not ; n3572
g3317 and b[29] b[30] ; n3573
g3318 and n3572_not n3573_not ; n3574
g3319 and n3571_not n3574 ; n3575
g3320 and n3571 n3574_not ; n3576
g3321 and n3575_not n3576_not ; n3577
g3322 and n269 n3577 ; n3578
g3323 and n3570 n3578_not ; n3579
g3324 and a[2] n3579_not ; n3580
g3325 and a[2] n3580_not ; n3581
g3326 and n3579_not n3580_not ; n3582
g3327 and n3581_not n3582_not ; n3583
g3328 and n3565 n3583_not ; n3584
g3329 and n3565 n3584_not ; n3585
g3330 and n3583_not n3584_not ; n3586
g3331 and n3585_not n3586_not ; n3587
g3332 and n3390_not n3395_not ; n3588
g3333 and n3587_not n3588_not ; n3589
g3334 and n3587 n3588 ; n3590
g3335 and n3589_not n3590_not ; f[30]
g3336 and b[16] n1302 ; n3592
g3337 and b[14] n1391 ; n3593
g3338 and b[15] n1297 ; n3594
g3339 and n3593_not n3594_not ; n3595
g3340 and n3592_not n3595 ; n3596
g3341 and n1237 n1305 ; n3597
g3342 and n3596 n3597_not ; n3598
g3343 and a[17] n3598_not ; n3599
g3344 and a[17] n3599_not ; n3600
g3345 and n3598_not n3599_not ; n3601
g3346 and n3600_not n3601_not ; n3602
g3347 and n3273_not n3458_not ; n3603
g3348 and n3455_not n3603_not ; n3604
g3349 and b[7] n2539 ; n3605
g3350 and b[5] n2685 ; n3606
g3351 and b[6] n2534 ; n3607
g3352 and n3606_not n3607_not ; n3608
g3353 and n3605_not n3608 ; n3609
g3354 and n484 n2542 ; n3610
g3355 and n3609 n3610_not ; n3611
g3356 and a[26] n3611_not ; n3612
g3357 and a[26] n3612_not ; n3613
g3358 and n3611_not n3612_not ; n3614
g3359 and n3613_not n3614_not ; n3615
g3360 and n3255 n3437 ; n3616
g3361 and n3452_not n3616_not ; n3617
g3362 and b[4] n3050 ; n3618
g3363 and b[2] n3243 ; n3619
g3364 and b[3] n3045 ; n3620
g3365 and n3619_not n3620_not ; n3621
g3366 and n3618_not n3621 ; n3622
g3367 and n346 n3053 ; n3623
g3368 and n3622 n3623_not ; n3624
g3369 and a[29] n3624_not ; n3625
g3370 and a[29] n3625_not ; n3626
g3371 and n3624_not n3625_not ; n3627
g3372 and n3626_not n3627_not ; n3628
g3373 and a[32] n3437_not ; n3629
g3374 and a[30]_not a[31] ; n3630
g3375 and a[30] a[31]_not ; n3631
g3376 and n3630_not n3631_not ; n3632
g3377 and n3436 n3632_not ; n3633
g3378 and b[0] n3633 ; n3634
g3379 and a[31]_not a[32] ; n3635
g3380 and a[31] a[32]_not ; n3636
g3381 and n3635_not n3636_not ; n3637
g3382 and n3436_not n3637 ; n3638
g3383 and b[1] n3638 ; n3639
g3384 and n3634_not n3639_not ; n3640
g3385 and n3436_not n3637_not ; n3641
g3386 and n272_not n3641 ; n3642
g3387 and n3640 n3642_not ; n3643
g3388 and a[32] n3643_not ; n3644
g3389 and a[32] n3644_not ; n3645
g3390 and n3643_not n3644_not ; n3646
g3391 and n3645_not n3646_not ; n3647
g3392 and n3629 n3647_not ; n3648
g3393 and n3629_not n3647 ; n3649
g3394 and n3648_not n3649_not ; n3650
g3395 and n3628 n3650 ; n3651
g3396 and n3628_not n3650_not ; n3652
g3397 and n3651_not n3652_not ; n3653
g3398 and n3617_not n3653_not ; n3654
g3399 and n3617 n3653 ; n3655
g3400 and n3654_not n3655_not ; n3656
g3401 and n3615_not n3656 ; n3657
g3402 and n3615 n3656_not ; n3658
g3403 and n3657_not n3658_not ; n3659
g3404 and n3604_not n3659 ; n3660
g3405 and n3604 n3659_not ; n3661
g3406 and n3660_not n3661_not ; n3662
g3407 and b[10] n2048 ; n3663
g3408 and b[8] n2198 ; n3664
g3409 and b[9] n2043 ; n3665
g3410 and n3664_not n3665_not ; n3666
g3411 and n3663_not n3666 ; n3667
g3412 and n738 n2051 ; n3668
g3413 and n3667 n3668_not ; n3669
g3414 and a[23] n3669_not ; n3670
g3415 and a[23] n3670_not ; n3671
g3416 and n3669_not n3670_not ; n3672
g3417 and n3671_not n3672_not ; n3673
g3418 and n3662 n3673_not ; n3674
g3419 and n3662 n3674_not ; n3675
g3420 and n3673_not n3674_not ; n3676
g3421 and n3675_not n3676_not ; n3677
g3422 and n3473_not n3476_not ; n3678
g3423 and n3677 n3678 ; n3679
g3424 and n3677_not n3678_not ; n3680
g3425 and n3679_not n3680_not ; n3681
g3426 and b[13] n1627 ; n3682
g3427 and b[11] n1763 ; n3683
g3428 and b[12] n1622 ; n3684
g3429 and n3683_not n3684_not ; n3685
g3430 and n3682_not n3685 ; n3686
g3431 and n1008 n1630 ; n3687
g3432 and n3686 n3687_not ; n3688
g3433 and a[20] n3688_not ; n3689
g3434 and a[20] n3689_not ; n3690
g3435 and n3688_not n3689_not ; n3691
g3436 and n3690_not n3691_not ; n3692
g3437 and n3681_not n3692 ; n3693
g3438 and n3681 n3692_not ; n3694
g3439 and n3693_not n3694_not ; n3695
g3440 and n3480_not n3482_not ; n3696
g3441 and n3695 n3696_not ; n3697
g3442 and n3695_not n3696 ; n3698
g3443 and n3697_not n3698_not ; n3699
g3444 and n3602_not n3699 ; n3700
g3445 and n3699 n3700_not ; n3701
g3446 and n3602_not n3700_not ; n3702
g3447 and n3701_not n3702_not ; n3703
g3448 and n3485_not n3491_not ; n3704
g3449 and n3703 n3704 ; n3705
g3450 and n3703_not n3704_not ; n3706
g3451 and n3705_not n3706_not ; n3707
g3452 and b[19] n951 ; n3708
g3453 and b[17] n1056 ; n3709
g3454 and b[18] n946 ; n3710
g3455 and n3709_not n3710_not ; n3711
g3456 and n3708_not n3711 ; n3712
g3457 and n954 n1708 ; n3713
g3458 and n3712 n3713_not ; n3714
g3459 and a[14] n3714_not ; n3715
g3460 and a[14] n3715_not ; n3716
g3461 and n3714_not n3715_not ; n3717
g3462 and n3716_not n3717_not ; n3718
g3463 and n3707 n3718_not ; n3719
g3464 and n3707 n3719_not ; n3720
g3465 and n3718_not n3719_not ; n3721
g3466 and n3720_not n3721_not ; n3722
g3467 and n3504_not n3510_not ; n3723
g3468 and n3722 n3723 ; n3724
g3469 and n3722_not n3723_not ; n3725
g3470 and n3724_not n3725_not ; n3726
g3471 and b[22] n700 ; n3727
g3472 and b[20] n767 ; n3728
g3473 and b[21] n695 ; n3729
g3474 and n3728_not n3729_not ; n3730
g3475 and n3727_not n3730 ; n3731
g3476 and n703 n2145 ; n3732
g3477 and n3731 n3732_not ; n3733
g3478 and a[11] n3733_not ; n3734
g3479 and a[11] n3734_not ; n3735
g3480 and n3733_not n3734_not ; n3736
g3481 and n3735_not n3736_not ; n3737
g3482 and n3726 n3737_not ; n3738
g3483 and n3726 n3738_not ; n3739
g3484 and n3737_not n3738_not ; n3740
g3485 and n3739_not n3740_not ; n3741
g3486 and n3342_not n3526_not ; n3742
g3487 and n3523_not n3742_not ; n3743
g3488 and n3741 n3743 ; n3744
g3489 and n3741_not n3743_not ; n3745
g3490 and n3744_not n3745_not ; n3746
g3491 and b[25] n511 ; n3747
g3492 and b[23] n541 ; n3748
g3493 and b[24] n506 ; n3749
g3494 and n3748_not n3749_not ; n3750
g3495 and n3747_not n3750 ; n3751
g3496 and n514 n2485 ; n3752
g3497 and n3751 n3752_not ; n3753
g3498 and a[8] n3753_not ; n3754
g3499 and a[8] n3754_not ; n3755
g3500 and n3753_not n3754_not ; n3756
g3501 and n3755_not n3756_not ; n3757
g3502 and n3746 n3757_not ; n3758
g3503 and n3746 n3758_not ; n3759
g3504 and n3757_not n3758_not ; n3760
g3505 and n3759_not n3760_not ; n3761
g3506 and n3541_not n3545_not ; n3762
g3507 and n3761 n3762 ; n3763
g3508 and n3761_not n3762_not ; n3764
g3509 and n3763_not n3764_not ; n3765
g3510 and b[28] n362 ; n3766
g3511 and b[26] n403 ; n3767
g3512 and b[27] n357 ; n3768
g3513 and n3767_not n3768_not ; n3769
g3514 and n3766_not n3769 ; n3770
g3515 and n365 n3189 ; n3771
g3516 and n3770 n3771_not ; n3772
g3517 and a[5] n3772_not ; n3773
g3518 and a[5] n3773_not ; n3774
g3519 and n3772_not n3773_not ; n3775
g3520 and n3774_not n3775_not ; n3776
g3521 and n3765 n3776_not ; n3777
g3522 and n3765 n3777_not ; n3778
g3523 and n3776_not n3777_not ; n3779
g3524 and n3778_not n3779_not ; n3780
g3525 and n3558_not n3564_not ; n3781
g3526 and n3780 n3781 ; n3782
g3527 and n3780_not n3781_not ; n3783
g3528 and n3782_not n3783_not ; n3784
g3529 and b[31] n266 ; n3785
g3530 and b[29] n284 ; n3786
g3531 and b[30] n261 ; n3787
g3532 and n3786_not n3787_not ; n3788
g3533 and n3785_not n3788 ; n3789
g3534 and n3573_not n3575_not ; n3790
g3535 and b[30]_not b[31]_not ; n3791
g3536 and b[30] b[31] ; n3792
g3537 and n3791_not n3792_not ; n3793
g3538 and n3790_not n3793 ; n3794
g3539 and n3790 n3793_not ; n3795
g3540 and n3794_not n3795_not ; n3796
g3541 and n269 n3796 ; n3797
g3542 and n3789 n3797_not ; n3798
g3543 and a[2] n3798_not ; n3799
g3544 and a[2] n3799_not ; n3800
g3545 and n3798_not n3799_not ; n3801
g3546 and n3800_not n3801_not ; n3802
g3547 and n3784 n3802_not ; n3803
g3548 and n3784 n3803_not ; n3804
g3549 and n3802_not n3803_not ; n3805
g3550 and n3804_not n3805_not ; n3806
g3551 and n3584_not n3589_not ; n3807
g3552 and n3806_not n3807_not ; n3808
g3553 and n3806 n3807 ; n3809
g3554 and n3808_not n3809_not ; f[31]
g3555 and n3803_not n3808_not ; n3811
g3556 and n3777_not n3783_not ; n3812
g3557 and b[26] n511 ; n3813
g3558 and b[24] n541 ; n3814
g3559 and b[25] n506 ; n3815
g3560 and n3814_not n3815_not ; n3816
g3561 and n3813_not n3816 ; n3817
g3562 and n514 n2813 ; n3818
g3563 and n3817 n3818_not ; n3819
g3564 and a[8] n3819_not ; n3820
g3565 and a[8] n3820_not ; n3821
g3566 and n3819_not n3820_not ; n3822
g3567 and n3821_not n3822_not ; n3823
g3568 and n3738_not n3745_not ; n3824
g3569 and n3719_not n3725_not ; n3825
g3570 and b[17] n1302 ; n3826
g3571 and b[15] n1391 ; n3827
g3572 and b[16] n1297 ; n3828
g3573 and n3827_not n3828_not ; n3829
g3574 and n3826_not n3829 ; n3830
g3575 and n1305 n1356 ; n3831
g3576 and n3830 n3831_not ; n3832
g3577 and a[17] n3832_not ; n3833
g3578 and a[17] n3833_not ; n3834
g3579 and n3832_not n3833_not ; n3835
g3580 and n3834_not n3835_not ; n3836
g3581 and n3694_not n3697_not ; n3837
g3582 and n3674_not n3680_not ; n3838
g3583 and n3628_not n3650 ; n3839
g3584 and n3654_not n3839_not ; n3840
g3585 and b[2] n3638 ; n3841
g3586 and n3436 n3637_not ; n3842
g3587 and n3632 n3842 ; n3843
g3588 and b[0] n3843 ; n3844
g3589 and b[1] n3633 ; n3845
g3590 and n3844_not n3845_not ; n3846
g3591 and n3841_not n3846 ; n3847
g3592 and n296 n3641 ; n3848
g3593 and n3847 n3848_not ; n3849
g3594 and a[32] n3849_not ; n3850
g3595 and a[32] n3850_not ; n3851
g3596 and n3849_not n3850_not ; n3852
g3597 and n3851_not n3852_not ; n3853
g3598 and n3648_not n3853 ; n3854
g3599 and n3648 n3853_not ; n3855
g3600 and n3854_not n3855_not ; n3856
g3601 and b[5] n3050 ; n3857
g3602 and b[3] n3243 ; n3858
g3603 and b[4] n3045 ; n3859
g3604 and n3858_not n3859_not ; n3860
g3605 and n3857_not n3860 ; n3861
g3606 and n394 n3053 ; n3862
g3607 and n3861 n3862_not ; n3863
g3608 and a[29] n3863_not ; n3864
g3609 and a[29] n3864_not ; n3865
g3610 and n3863_not n3864_not ; n3866
g3611 and n3865_not n3866_not ; n3867
g3612 and n3856 n3867_not ; n3868
g3613 and n3856_not n3867 ; n3869
g3614 and n3840_not n3869_not ; n3870
g3615 and n3868_not n3870 ; n3871
g3616 and n3840_not n3871_not ; n3872
g3617 and n3868_not n3871_not ; n3873
g3618 and n3869_not n3873 ; n3874
g3619 and n3872_not n3874_not ; n3875
g3620 and b[8] n2539 ; n3876
g3621 and b[6] n2685 ; n3877
g3622 and b[7] n2534 ; n3878
g3623 and n3877_not n3878_not ; n3879
g3624 and n3876_not n3879 ; n3880
g3625 and n585 n2542 ; n3881
g3626 and n3880 n3881_not ; n3882
g3627 and a[26] n3882_not ; n3883
g3628 and a[26] n3883_not ; n3884
g3629 and n3882_not n3883_not ; n3885
g3630 and n3884_not n3885_not ; n3886
g3631 and n3875_not n3886_not ; n3887
g3632 and n3875_not n3887_not ; n3888
g3633 and n3886_not n3887_not ; n3889
g3634 and n3888_not n3889_not ; n3890
g3635 and n3657_not n3660_not ; n3891
g3636 and n3890 n3891 ; n3892
g3637 and n3890_not n3891_not ; n3893
g3638 and n3892_not n3893_not ; n3894
g3639 and b[11] n2048 ; n3895
g3640 and b[9] n2198 ; n3896
g3641 and b[10] n2043 ; n3897
g3642 and n3896_not n3897_not ; n3898
g3643 and n3895_not n3898 ; n3899
g3644 and n818 n2051 ; n3900
g3645 and n3899 n3900_not ; n3901
g3646 and a[23] n3901_not ; n3902
g3647 and a[23] n3902_not ; n3903
g3648 and n3901_not n3902_not ; n3904
g3649 and n3903_not n3904_not ; n3905
g3650 and n3894 n3905_not ; n3906
g3651 and n3894_not n3905 ; n3907
g3652 and n3838_not n3907_not ; n3908
g3653 and n3906_not n3908 ; n3909
g3654 and n3838_not n3909_not ; n3910
g3655 and n3906_not n3909_not ; n3911
g3656 and n3907_not n3911 ; n3912
g3657 and n3910_not n3912_not ; n3913
g3658 and b[14] n1627 ; n3914
g3659 and b[12] n1763 ; n3915
g3660 and b[13] n1622 ; n3916
g3661 and n3915_not n3916_not ; n3917
g3662 and n3914_not n3917 ; n3918
g3663 and n1034 n1630 ; n3919
g3664 and n3918 n3919_not ; n3920
g3665 and a[20] n3920_not ; n3921
g3666 and a[20] n3921_not ; n3922
g3667 and n3920_not n3921_not ; n3923
g3668 and n3922_not n3923_not ; n3924
g3669 and n3913 n3924 ; n3925
g3670 and n3913_not n3924_not ; n3926
g3671 and n3925_not n3926_not ; n3927
g3672 and n3837_not n3927 ; n3928
g3673 and n3837 n3927_not ; n3929
g3674 and n3928_not n3929_not ; n3930
g3675 and n3836_not n3930 ; n3931
g3676 and n3930 n3931_not ; n3932
g3677 and n3836_not n3931_not ; n3933
g3678 and n3932_not n3933_not ; n3934
g3679 and n3700_not n3706_not ; n3935
g3680 and n3934 n3935 ; n3936
g3681 and n3934_not n3935_not ; n3937
g3682 and n3936_not n3937_not ; n3938
g3683 and b[20] n951 ; n3939
g3684 and b[18] n1056 ; n3940
g3685 and b[19] n946 ; n3941
g3686 and n3940_not n3941_not ; n3942
g3687 and n3939_not n3942 ; n3943
g3688 and n954 n1846 ; n3944
g3689 and n3943 n3944_not ; n3945
g3690 and a[14] n3945_not ; n3946
g3691 and a[14] n3946_not ; n3947
g3692 and n3945_not n3946_not ; n3948
g3693 and n3947_not n3948_not ; n3949
g3694 and n3938 n3949_not ; n3950
g3695 and n3938_not n3949 ; n3951
g3696 and n3825_not n3951_not ; n3952
g3697 and n3950_not n3952 ; n3953
g3698 and n3825_not n3953_not ; n3954
g3699 and n3950_not n3953_not ; n3955
g3700 and n3951_not n3955 ; n3956
g3701 and n3954_not n3956_not ; n3957
g3702 and b[23] n700 ; n3958
g3703 and b[21] n767 ; n3959
g3704 and b[22] n695 ; n3960
g3705 and n3959_not n3960_not ; n3961
g3706 and n3958_not n3961 ; n3962
g3707 and n703 n2300 ; n3963
g3708 and n3962 n3963_not ; n3964
g3709 and a[11] n3964_not ; n3965
g3710 and a[11] n3965_not ; n3966
g3711 and n3964_not n3965_not ; n3967
g3712 and n3966_not n3967_not ; n3968
g3713 and n3957 n3968 ; n3969
g3714 and n3957_not n3968_not ; n3970
g3715 and n3969_not n3970_not ; n3971
g3716 and n3824_not n3971 ; n3972
g3717 and n3824 n3971_not ; n3973
g3718 and n3972_not n3973_not ; n3974
g3719 and n3823_not n3974 ; n3975
g3720 and n3974 n3975_not ; n3976
g3721 and n3823_not n3975_not ; n3977
g3722 and n3976_not n3977_not ; n3978
g3723 and n3758_not n3764_not ; n3979
g3724 and n3978 n3979 ; n3980
g3725 and n3978_not n3979_not ; n3981
g3726 and n3980_not n3981_not ; n3982
g3727 and b[29] n362 ; n3983
g3728 and b[27] n403 ; n3984
g3729 and b[28] n357 ; n3985
g3730 and n3984_not n3985_not ; n3986
g3731 and n3983_not n3986 ; n3987
g3732 and n365 n3383 ; n3988
g3733 and n3987 n3988_not ; n3989
g3734 and a[5] n3989_not ; n3990
g3735 and a[5] n3990_not ; n3991
g3736 and n3989_not n3990_not ; n3992
g3737 and n3991_not n3992_not ; n3993
g3738 and n3982 n3993_not ; n3994
g3739 and n3982_not n3993 ; n3995
g3740 and n3812_not n3995_not ; n3996
g3741 and n3994_not n3996 ; n3997
g3742 and n3812_not n3997_not ; n3998
g3743 and n3994_not n3997_not ; n3999
g3744 and n3995_not n3999 ; n4000
g3745 and n3998_not n4000_not ; n4001
g3746 and b[32] n266 ; n4002
g3747 and b[30] n284 ; n4003
g3748 and b[31] n261 ; n4004
g3749 and n4003_not n4004_not ; n4005
g3750 and n4002_not n4005 ; n4006
g3751 and n3792_not n3794_not ; n4007
g3752 and b[31]_not b[32]_not ; n4008
g3753 and b[31] b[32] ; n4009
g3754 and n4008_not n4009_not ; n4010
g3755 and n4007_not n4010 ; n4011
g3756 and n4007 n4010_not ; n4012
g3757 and n4011_not n4012_not ; n4013
g3758 and n269 n4013 ; n4014
g3759 and n4006 n4014_not ; n4015
g3760 and a[2] n4015_not ; n4016
g3761 and a[2] n4016_not ; n4017
g3762 and n4015_not n4016_not ; n4018
g3763 and n4017_not n4018_not ; n4019
g3764 and n4001_not n4019 ; n4020
g3765 and n4001 n4019_not ; n4021
g3766 and n4020_not n4021_not ; n4022
g3767 and n3811_not n4022_not ; n4023
g3768 and n3811 n4022 ; n4024
g3769 and n4023_not n4024_not ; f[32]
g3770 and n4001_not n4019_not ; n4026
g3771 and n4023_not n4026_not ; n4027
g3772 and b[27] n511 ; n4028
g3773 and b[25] n541 ; n4029
g3774 and b[26] n506 ; n4030
g3775 and n4029_not n4030_not ; n4031
g3776 and n4028_not n4031 ; n4032
g3777 and n514 n2990 ; n4033
g3778 and n4032 n4033_not ; n4034
g3779 and a[8] n4034_not ; n4035
g3780 and a[8] n4035_not ; n4036
g3781 and n4034_not n4035_not ; n4037
g3782 and n4036_not n4037_not ; n4038
g3783 and n3970_not n3972_not ; n4039
g3784 and n3931_not n3937_not ; n4040
g3785 and n3926_not n3928_not ; n4041
g3786 and b[15] n1627 ; n4042
g3787 and b[13] n1763 ; n4043
g3788 and b[14] n1622 ; n4044
g3789 and n4043_not n4044_not ; n4045
g3790 and n4042_not n4045 ; n4046
g3791 and n1131 n1630 ; n4047
g3792 and n4046 n4047_not ; n4048
g3793 and a[20] n4048_not ; n4049
g3794 and a[20] n4049_not ; n4050
g3795 and n4048_not n4049_not ; n4051
g3796 and n4050_not n4051_not ; n4052
g3797 and n3887_not n3893_not ; n4053
g3798 and b[6] n3050 ; n4054
g3799 and b[4] n3243 ; n4055
g3800 and b[5] n3045 ; n4056
g3801 and n4055_not n4056_not ; n4057
g3802 and n4054_not n4057 ; n4058
g3803 and n459 n3053 ; n4059
g3804 and n4058 n4059_not ; n4060
g3805 and a[29] n4060_not ; n4061
g3806 and a[29] n4061_not ; n4062
g3807 and n4060_not n4061_not ; n4063
g3808 and n4062_not n4063_not ; n4064
g3809 and a[32] a[33]_not ; n4065
g3810 and a[32]_not a[33] ; n4066
g3811 and n4065_not n4066_not ; n4067
g3812 and b[0] n4067_not ; n4068
g3813 and n3855_not n4068 ; n4069
g3814 and n3855 n4068_not ; n4070
g3815 and n4069_not n4070_not ; n4071
g3816 and b[3] n3638 ; n4072
g3817 and b[1] n3843 ; n4073
g3818 and b[2] n3633 ; n4074
g3819 and n4073_not n4074_not ; n4075
g3820 and n4072_not n4075 ; n4076
g3821 and n318 n3641 ; n4077
g3822 and n4076 n4077_not ; n4078
g3823 and a[32] n4078_not ; n4079
g3824 and a[32] n4079_not ; n4080
g3825 and n4078_not n4079_not ; n4081
g3826 and n4080_not n4081_not ; n4082
g3827 and n4071_not n4082_not ; n4083
g3828 and n4071 n4082 ; n4084
g3829 and n4083_not n4084_not ; n4085
g3830 and n4064_not n4085 ; n4086
g3831 and n4085 n4086_not ; n4087
g3832 and n4064_not n4086_not ; n4088
g3833 and n4087_not n4088_not ; n4089
g3834 and n3873_not n4089 ; n4090
g3835 and n3873 n4089_not ; n4091
g3836 and n4090_not n4091_not ; n4092
g3837 and b[9] n2539 ; n4093
g3838 and b[7] n2685 ; n4094
g3839 and b[8] n2534 ; n4095
g3840 and n4094_not n4095_not ; n4096
g3841 and n4093_not n4096 ; n4097
g3842 and n651 n2542 ; n4098
g3843 and n4097 n4098_not ; n4099
g3844 and a[26] n4099_not ; n4100
g3845 and a[26] n4100_not ; n4101
g3846 and n4099_not n4100_not ; n4102
g3847 and n4101_not n4102_not ; n4103
g3848 and n4092_not n4103_not ; n4104
g3849 and n4092 n4103 ; n4105
g3850 and n4104_not n4105_not ; n4106
g3851 and n4053 n4106_not ; n4107
g3852 and n4053_not n4106 ; n4108
g3853 and n4107_not n4108_not ; n4109
g3854 and b[12] n2048 ; n4110
g3855 and b[10] n2198 ; n4111
g3856 and b[11] n2043 ; n4112
g3857 and n4111_not n4112_not ; n4113
g3858 and n4110_not n4113 ; n4114
g3859 and n842 n2051 ; n4115
g3860 and n4114 n4115_not ; n4116
g3861 and a[23] n4116_not ; n4117
g3862 and a[23] n4117_not ; n4118
g3863 and n4116_not n4117_not ; n4119
g3864 and n4118_not n4119_not ; n4120
g3865 and n4109_not n4120 ; n4121
g3866 and n4109 n4120_not ; n4122
g3867 and n4121_not n4122_not ; n4123
g3868 and n3911_not n4123 ; n4124
g3869 and n3911 n4123_not ; n4125
g3870 and n4124_not n4125_not ; n4126
g3871 and n4052_not n4126 ; n4127
g3872 and n4126 n4127_not ; n4128
g3873 and n4052_not n4127_not ; n4129
g3874 and n4128_not n4129_not ; n4130
g3875 and n4041_not n4130 ; n4131
g3876 and n4041 n4130_not ; n4132
g3877 and n4131_not n4132_not ; n4133
g3878 and b[18] n1302 ; n4134
g3879 and b[16] n1391 ; n4135
g3880 and b[17] n1297 ; n4136
g3881 and n4135_not n4136_not ; n4137
g3882 and n4134_not n4137 ; n4138
g3883 and n1305 n1566 ; n4139
g3884 and n4138 n4139_not ; n4140
g3885 and a[17] n4140_not ; n4141
g3886 and a[17] n4141_not ; n4142
g3887 and n4140_not n4141_not ; n4143
g3888 and n4142_not n4143_not ; n4144
g3889 and n4133_not n4144_not ; n4145
g3890 and n4133 n4144 ; n4146
g3891 and n4145_not n4146_not ; n4147
g3892 and n4040 n4147_not ; n4148
g3893 and n4040_not n4147 ; n4149
g3894 and n4148_not n4149_not ; n4150
g3895 and b[21] n951 ; n4151
g3896 and b[19] n1056 ; n4152
g3897 and b[20] n946 ; n4153
g3898 and n4152_not n4153_not ; n4154
g3899 and n4151_not n4154 ; n4155
g3900 and n954 n1984 ; n4156
g3901 and n4155 n4156_not ; n4157
g3902 and a[14] n4157_not ; n4158
g3903 and a[14] n4158_not ; n4159
g3904 and n4157_not n4158_not ; n4160
g3905 and n4159_not n4160_not ; n4161
g3906 and n4150 n4161_not ; n4162
g3907 and n4150 n4162_not ; n4163
g3908 and n4161_not n4162_not ; n4164
g3909 and n4163_not n4164_not ; n4165
g3910 and n3955_not n4165 ; n4166
g3911 and n3955 n4165_not ; n4167
g3912 and n4166_not n4167_not ; n4168
g3913 and b[24] n700 ; n4169
g3914 and b[22] n767 ; n4170
g3915 and b[23] n695 ; n4171
g3916 and n4170_not n4171_not ; n4172
g3917 and n4169_not n4172 ; n4173
g3918 and n703 n2458 ; n4174
g3919 and n4173 n4174_not ; n4175
g3920 and a[11] n4175_not ; n4176
g3921 and a[11] n4176_not ; n4177
g3922 and n4175_not n4176_not ; n4178
g3923 and n4177_not n4178_not ; n4179
g3924 and n4168 n4179 ; n4180
g3925 and n4168_not n4179_not ; n4181
g3926 and n4180_not n4181_not ; n4182
g3927 and n4039_not n4182 ; n4183
g3928 and n4039 n4182_not ; n4184
g3929 and n4183_not n4184_not ; n4185
g3930 and n4038_not n4185 ; n4186
g3931 and n4185 n4186_not ; n4187
g3932 and n4038_not n4186_not ; n4188
g3933 and n4187_not n4188_not ; n4189
g3934 and n3975_not n3981_not ; n4190
g3935 and n4189 n4190 ; n4191
g3936 and n4189_not n4190_not ; n4192
g3937 and n4191_not n4192_not ; n4193
g3938 and b[30] n362 ; n4194
g3939 and b[28] n403 ; n4195
g3940 and b[29] n357 ; n4196
g3941 and n4195_not n4196_not ; n4197
g3942 and n4194_not n4197 ; n4198
g3943 and n365 n3577 ; n4199
g3944 and n4198 n4199_not ; n4200
g3945 and a[5] n4200_not ; n4201
g3946 and a[5] n4201_not ; n4202
g3947 and n4200_not n4201_not ; n4203
g3948 and n4202_not n4203_not ; n4204
g3949 and n4193 n4204_not ; n4205
g3950 and n4193 n4205_not ; n4206
g3951 and n4204_not n4205_not ; n4207
g3952 and n4206_not n4207_not ; n4208
g3953 and n3999_not n4208 ; n4209
g3954 and n3999 n4208_not ; n4210
g3955 and n4209_not n4210_not ; n4211
g3956 and b[33] n266 ; n4212
g3957 and b[31] n284 ; n4213
g3958 and b[32] n261 ; n4214
g3959 and n4213_not n4214_not ; n4215
g3960 and n4212_not n4215 ; n4216
g3961 and n4009_not n4011_not ; n4217
g3962 and b[32]_not b[33]_not ; n4218
g3963 and b[32] b[33] ; n4219
g3964 and n4218_not n4219_not ; n4220
g3965 and n4217_not n4220 ; n4221
g3966 and n4217 n4220_not ; n4222
g3967 and n4221_not n4222_not ; n4223
g3968 and n269 n4223 ; n4224
g3969 and n4216 n4224_not ; n4225
g3970 and a[2] n4225_not ; n4226
g3971 and a[2] n4226_not ; n4227
g3972 and n4225_not n4226_not ; n4228
g3973 and n4227_not n4228_not ; n4229
g3974 and n4211_not n4229_not ; n4230
g3975 and n4211 n4229 ; n4231
g3976 and n4230_not n4231_not ; n4232
g3977 and n4027_not n4232 ; n4233
g3978 and n4027 n4232_not ; n4234
g3979 and n4233_not n4234_not ; f[33]
g3980 and n4230_not n4233_not ; n4236
g3981 and n3999_not n4208_not ; n4237
g3982 and n4205_not n4237_not ; n4238
g3983 and n4181_not n4183_not ; n4239
g3984 and n4122_not n4124_not ; n4240
g3985 and b[10] n2539 ; n4241
g3986 and b[8] n2685 ; n4242
g3987 and b[9] n2534 ; n4243
g3988 and n4242_not n4243_not ; n4244
g3989 and n4241_not n4244 ; n4245
g3990 and n738 n2542 ; n4246
g3991 and n4245 n4246_not ; n4247
g3992 and a[26] n4247_not ; n4248
g3993 and a[26] n4248_not ; n4249
g3994 and n4247_not n4248_not ; n4250
g3995 and n4249_not n4250_not ; n4251
g3996 and n3873_not n4089_not ; n4252
g3997 and n4086_not n4252_not ; n4253
g3998 and b[7] n3050 ; n4254
g3999 and b[5] n3243 ; n4255
g4000 and b[6] n3045 ; n4256
g4001 and n4255_not n4256_not ; n4257
g4002 and n4254_not n4257 ; n4258
g4003 and n484 n3053 ; n4259
g4004 and n4258 n4259_not ; n4260
g4005 and a[29] n4260_not ; n4261
g4006 and a[29] n4261_not ; n4262
g4007 and n4260_not n4261_not ; n4263
g4008 and n4262_not n4263_not ; n4264
g4009 and n3855 n4068 ; n4265
g4010 and n4083_not n4265_not ; n4266
g4011 and b[4] n3638 ; n4267
g4012 and b[2] n3843 ; n4268
g4013 and b[3] n3633 ; n4269
g4014 and n4268_not n4269_not ; n4270
g4015 and n4267_not n4270 ; n4271
g4016 and n346 n3641 ; n4272
g4017 and n4271 n4272_not ; n4273
g4018 and a[32] n4273_not ; n4274
g4019 and a[32] n4274_not ; n4275
g4020 and n4273_not n4274_not ; n4276
g4021 and n4275_not n4276_not ; n4277
g4022 and a[35] n4068_not ; n4278
g4023 and a[33]_not a[34] ; n4279
g4024 and a[33] a[34]_not ; n4280
g4025 and n4279_not n4280_not ; n4281
g4026 and n4067 n4281_not ; n4282
g4027 and b[0] n4282 ; n4283
g4028 and a[34]_not a[35] ; n4284
g4029 and a[34] a[35]_not ; n4285
g4030 and n4284_not n4285_not ; n4286
g4031 and n4067_not n4286 ; n4287
g4032 and b[1] n4287 ; n4288
g4033 and n4283_not n4288_not ; n4289
g4034 and n4067_not n4286_not ; n4290
g4035 and n272_not n4290 ; n4291
g4036 and n4289 n4291_not ; n4292
g4037 and a[35] n4292_not ; n4293
g4038 and a[35] n4293_not ; n4294
g4039 and n4292_not n4293_not ; n4295
g4040 and n4294_not n4295_not ; n4296
g4041 and n4278 n4296_not ; n4297
g4042 and n4278_not n4296 ; n4298
g4043 and n4297_not n4298_not ; n4299
g4044 and n4277 n4299_not ; n4300
g4045 and n4277_not n4299 ; n4301
g4046 and n4300_not n4301_not ; n4302
g4047 and n4266_not n4302 ; n4303
g4048 and n4266 n4302_not ; n4304
g4049 and n4303_not n4304_not ; n4305
g4050 and n4264 n4305_not ; n4306
g4051 and n4264_not n4305 ; n4307
g4052 and n4306_not n4307_not ; n4308
g4053 and n4253_not n4308 ; n4309
g4054 and n4253 n4308_not ; n4310
g4055 and n4309_not n4310_not ; n4311
g4056 and n4251_not n4311 ; n4312
g4057 and n4311 n4312_not ; n4313
g4058 and n4251_not n4312_not ; n4314
g4059 and n4313_not n4314_not ; n4315
g4060 and n4104_not n4108_not ; n4316
g4061 and n4315 n4316 ; n4317
g4062 and n4315_not n4316_not ; n4318
g4063 and n4317_not n4318_not ; n4319
g4064 and b[13] n2048 ; n4320
g4065 and b[11] n2198 ; n4321
g4066 and b[12] n2043 ; n4322
g4067 and n4321_not n4322_not ; n4323
g4068 and n4320_not n4323 ; n4324
g4069 and n1008 n2051 ; n4325
g4070 and n4324 n4325_not ; n4326
g4071 and a[23] n4326_not ; n4327
g4072 and a[23] n4327_not ; n4328
g4073 and n4326_not n4327_not ; n4329
g4074 and n4328_not n4329_not ; n4330
g4075 and n4319 n4330_not ; n4331
g4076 and n4319_not n4330 ; n4332
g4077 and n4240_not n4332_not ; n4333
g4078 and n4331_not n4333 ; n4334
g4079 and n4240_not n4334_not ; n4335
g4080 and n4331_not n4334_not ; n4336
g4081 and n4332_not n4336 ; n4337
g4082 and n4335_not n4337_not ; n4338
g4083 and b[16] n1627 ; n4339
g4084 and b[14] n1763 ; n4340
g4085 and b[15] n1622 ; n4341
g4086 and n4340_not n4341_not ; n4342
g4087 and n4339_not n4342 ; n4343
g4088 and n1237 n1630 ; n4344
g4089 and n4343 n4344_not ; n4345
g4090 and a[20] n4345_not ; n4346
g4091 and a[20] n4346_not ; n4347
g4092 and n4345_not n4346_not ; n4348
g4093 and n4347_not n4348_not ; n4349
g4094 and n4338_not n4349_not ; n4350
g4095 and n4338_not n4350_not ; n4351
g4096 and n4349_not n4350_not ; n4352
g4097 and n4351_not n4352_not ; n4353
g4098 and n4041_not n4130_not ; n4354
g4099 and n4127_not n4354_not ; n4355
g4100 and n4353 n4355 ; n4356
g4101 and n4353_not n4355_not ; n4357
g4102 and n4356_not n4357_not ; n4358
g4103 and b[19] n1302 ; n4359
g4104 and b[17] n1391 ; n4360
g4105 and b[18] n1297 ; n4361
g4106 and n4360_not n4361_not ; n4362
g4107 and n4359_not n4362 ; n4363
g4108 and n1305 n1708 ; n4364
g4109 and n4363 n4364_not ; n4365
g4110 and a[17] n4365_not ; n4366
g4111 and a[17] n4366_not ; n4367
g4112 and n4365_not n4366_not ; n4368
g4113 and n4367_not n4368_not ; n4369
g4114 and n4358 n4369_not ; n4370
g4115 and n4358 n4370_not ; n4371
g4116 and n4369_not n4370_not ; n4372
g4117 and n4371_not n4372_not ; n4373
g4118 and n4145_not n4149_not ; n4374
g4119 and n4373 n4374 ; n4375
g4120 and n4373_not n4374_not ; n4376
g4121 and n4375_not n4376_not ; n4377
g4122 and b[22] n951 ; n4378
g4123 and b[20] n1056 ; n4379
g4124 and b[21] n946 ; n4380
g4125 and n4379_not n4380_not ; n4381
g4126 and n4378_not n4381 ; n4382
g4127 and n954 n2145 ; n4383
g4128 and n4382 n4383_not ; n4384
g4129 and a[14] n4384_not ; n4385
g4130 and a[14] n4385_not ; n4386
g4131 and n4384_not n4385_not ; n4387
g4132 and n4386_not n4387_not ; n4388
g4133 and n4377 n4388_not ; n4389
g4134 and n4377 n4389_not ; n4390
g4135 and n4388_not n4389_not ; n4391
g4136 and n4390_not n4391_not ; n4392
g4137 and n3955_not n4165_not ; n4393
g4138 and n4162_not n4393_not ; n4394
g4139 and n4392 n4394 ; n4395
g4140 and n4392_not n4394_not ; n4396
g4141 and n4395_not n4396_not ; n4397
g4142 and b[25] n700 ; n4398
g4143 and b[23] n767 ; n4399
g4144 and b[24] n695 ; n4400
g4145 and n4399_not n4400_not ; n4401
g4146 and n4398_not n4401 ; n4402
g4147 and n703 n2485 ; n4403
g4148 and n4402 n4403_not ; n4404
g4149 and a[11] n4404_not ; n4405
g4150 and a[11] n4405_not ; n4406
g4151 and n4404_not n4405_not ; n4407
g4152 and n4406_not n4407_not ; n4408
g4153 and n4397 n4408_not ; n4409
g4154 and n4397_not n4408 ; n4410
g4155 and n4239_not n4410_not ; n4411
g4156 and n4409_not n4411 ; n4412
g4157 and n4239_not n4412_not ; n4413
g4158 and n4409_not n4412_not ; n4414
g4159 and n4410_not n4414 ; n4415
g4160 and n4413_not n4415_not ; n4416
g4161 and b[28] n511 ; n4417
g4162 and b[26] n541 ; n4418
g4163 and b[27] n506 ; n4419
g4164 and n4418_not n4419_not ; n4420
g4165 and n4417_not n4420 ; n4421
g4166 and n514 n3189 ; n4422
g4167 and n4421 n4422_not ; n4423
g4168 and a[8] n4423_not ; n4424
g4169 and a[8] n4424_not ; n4425
g4170 and n4423_not n4424_not ; n4426
g4171 and n4425_not n4426_not ; n4427
g4172 and n4416_not n4427_not ; n4428
g4173 and n4416_not n4428_not ; n4429
g4174 and n4427_not n4428_not ; n4430
g4175 and n4429_not n4430_not ; n4431
g4176 and n4186_not n4192_not ; n4432
g4177 and n4431 n4432 ; n4433
g4178 and n4431_not n4432_not ; n4434
g4179 and n4433_not n4434_not ; n4435
g4180 and b[31] n362 ; n4436
g4181 and b[29] n403 ; n4437
g4182 and b[30] n357 ; n4438
g4183 and n4437_not n4438_not ; n4439
g4184 and n4436_not n4439 ; n4440
g4185 and n365 n3796 ; n4441
g4186 and n4440 n4441_not ; n4442
g4187 and a[5] n4442_not ; n4443
g4188 and a[5] n4443_not ; n4444
g4189 and n4442_not n4443_not ; n4445
g4190 and n4444_not n4445_not ; n4446
g4191 and n4435 n4446_not ; n4447
g4192 and n4435_not n4446 ; n4448
g4193 and n4238_not n4448_not ; n4449
g4194 and n4447_not n4449 ; n4450
g4195 and n4238_not n4450_not ; n4451
g4196 and n4447_not n4450_not ; n4452
g4197 and n4448_not n4452 ; n4453
g4198 and n4451_not n4453_not ; n4454
g4199 and b[34] n266 ; n4455
g4200 and b[32] n284 ; n4456
g4201 and b[33] n261 ; n4457
g4202 and n4456_not n4457_not ; n4458
g4203 and n4455_not n4458 ; n4459
g4204 and n4219_not n4221_not ; n4460
g4205 and b[33]_not b[34]_not ; n4461
g4206 and b[33] b[34] ; n4462
g4207 and n4461_not n4462_not ; n4463
g4208 and n4460_not n4463 ; n4464
g4209 and n4460 n4463_not ; n4465
g4210 and n4464_not n4465_not ; n4466
g4211 and n269 n4466 ; n4467
g4212 and n4459 n4467_not ; n4468
g4213 and a[2] n4468_not ; n4469
g4214 and a[2] n4469_not ; n4470
g4215 and n4468_not n4469_not ; n4471
g4216 and n4470_not n4471_not ; n4472
g4217 and n4454_not n4472 ; n4473
g4218 and n4454 n4472_not ; n4474
g4219 and n4473_not n4474_not ; n4475
g4220 and n4236_not n4475_not ; n4476
g4221 and n4236 n4475 ; n4477
g4222 and n4476_not n4477_not ; f[34]
g4223 and n4454_not n4472_not ; n4479
g4224 and n4476_not n4479_not ; n4480
g4225 and b[29] n511 ; n4481
g4226 and b[27] n541 ; n4482
g4227 and b[28] n506 ; n4483
g4228 and n4482_not n4483_not ; n4484
g4229 and n4481_not n4484 ; n4485
g4230 and n514 n3383 ; n4486
g4231 and n4485 n4486_not ; n4487
g4232 and a[8] n4487_not ; n4488
g4233 and a[8] n4488_not ; n4489
g4234 and n4487_not n4488_not ; n4490
g4235 and n4489_not n4490_not ; n4491
g4236 and b[26] n700 ; n4492
g4237 and b[24] n767 ; n4493
g4238 and b[25] n695 ; n4494
g4239 and n4493_not n4494_not ; n4495
g4240 and n4492_not n4495 ; n4496
g4241 and n703 n2813 ; n4497
g4242 and n4496 n4497_not ; n4498
g4243 and a[11] n4498_not ; n4499
g4244 and a[11] n4499_not ; n4500
g4245 and n4498_not n4499_not ; n4501
g4246 and n4500_not n4501_not ; n4502
g4247 and n4389_not n4396_not ; n4503
g4248 and n4370_not n4376_not ; n4504
g4249 and b[17] n1627 ; n4505
g4250 and b[15] n1763 ; n4506
g4251 and b[16] n1622 ; n4507
g4252 and n4506_not n4507_not ; n4508
g4253 and n4505_not n4508 ; n4509
g4254 and n1356 n1630 ; n4510
g4255 and n4509 n4510_not ; n4511
g4256 and a[20] n4511_not ; n4512
g4257 and a[20] n4512_not ; n4513
g4258 and n4511_not n4512_not ; n4514
g4259 and n4513_not n4514_not ; n4515
g4260 and n4312_not n4318_not ; n4516
g4261 and b[11] n2539 ; n4517
g4262 and b[9] n2685 ; n4518
g4263 and b[10] n2534 ; n4519
g4264 and n4518_not n4519_not ; n4520
g4265 and n4517_not n4520 ; n4521
g4266 and n818 n2542 ; n4522
g4267 and n4521 n4522_not ; n4523
g4268 and a[26] n4523_not ; n4524
g4269 and a[26] n4524_not ; n4525
g4270 and n4523_not n4524_not ; n4526
g4271 and n4525_not n4526_not ; n4527
g4272 and n4307_not n4309_not ; n4528
g4273 and n4301_not n4303_not ; n4529
g4274 and b[2] n4287 ; n4530
g4275 and n4067 n4286_not ; n4531
g4276 and n4281 n4531 ; n4532
g4277 and b[0] n4532 ; n4533
g4278 and b[1] n4282 ; n4534
g4279 and n4533_not n4534_not ; n4535
g4280 and n4530_not n4535 ; n4536
g4281 and n296 n4290 ; n4537
g4282 and n4536 n4537_not ; n4538
g4283 and a[35] n4538_not ; n4539
g4284 and a[35] n4539_not ; n4540
g4285 and n4538_not n4539_not ; n4541
g4286 and n4540_not n4541_not ; n4542
g4287 and n4297_not n4542 ; n4543
g4288 and n4297 n4542_not ; n4544
g4289 and n4543_not n4544_not ; n4545
g4290 and b[5] n3638 ; n4546
g4291 and b[3] n3843 ; n4547
g4292 and b[4] n3633 ; n4548
g4293 and n4547_not n4548_not ; n4549
g4294 and n4546_not n4549 ; n4550
g4295 and n394 n3641 ; n4551
g4296 and n4550 n4551_not ; n4552
g4297 and a[32] n4552_not ; n4553
g4298 and a[32] n4553_not ; n4554
g4299 and n4552_not n4553_not ; n4555
g4300 and n4554_not n4555_not ; n4556
g4301 and n4545 n4556_not ; n4557
g4302 and n4545_not n4556 ; n4558
g4303 and n4529_not n4558_not ; n4559
g4304 and n4557_not n4559 ; n4560
g4305 and n4529_not n4560_not ; n4561
g4306 and n4557_not n4560_not ; n4562
g4307 and n4558_not n4562 ; n4563
g4308 and n4561_not n4563_not ; n4564
g4309 and b[8] n3050 ; n4565
g4310 and b[6] n3243 ; n4566
g4311 and b[7] n3045 ; n4567
g4312 and n4566_not n4567_not ; n4568
g4313 and n4565_not n4568 ; n4569
g4314 and n585 n3053 ; n4570
g4315 and n4569 n4570_not ; n4571
g4316 and a[29] n4571_not ; n4572
g4317 and a[29] n4572_not ; n4573
g4318 and n4571_not n4572_not ; n4574
g4319 and n4573_not n4574_not ; n4575
g4320 and n4564_not n4575_not ; n4576
g4321 and n4564_not n4576_not ; n4577
g4322 and n4575_not n4576_not ; n4578
g4323 and n4577_not n4578_not ; n4579
g4324 and n4528_not n4579_not ; n4580
g4325 and n4528 n4579 ; n4581
g4326 and n4580_not n4581_not ; n4582
g4327 and n4527_not n4582 ; n4583
g4328 and n4527_not n4583_not ; n4584
g4329 and n4582 n4583_not ; n4585
g4330 and n4584_not n4585_not ; n4586
g4331 and n4516_not n4586_not ; n4587
g4332 and n4516_not n4587_not ; n4588
g4333 and n4586_not n4587_not ; n4589
g4334 and n4588_not n4589_not ; n4590
g4335 and b[14] n2048 ; n4591
g4336 and b[12] n2198 ; n4592
g4337 and b[13] n2043 ; n4593
g4338 and n4592_not n4593_not ; n4594
g4339 and n4591_not n4594 ; n4595
g4340 and n1034 n2051 ; n4596
g4341 and n4595 n4596_not ; n4597
g4342 and a[23] n4597_not ; n4598
g4343 and a[23] n4598_not ; n4599
g4344 and n4597_not n4598_not ; n4600
g4345 and n4599_not n4600_not ; n4601
g4346 and n4590 n4601 ; n4602
g4347 and n4590_not n4601_not ; n4603
g4348 and n4602_not n4603_not ; n4604
g4349 and n4336_not n4604 ; n4605
g4350 and n4336 n4604_not ; n4606
g4351 and n4605_not n4606_not ; n4607
g4352 and n4515_not n4607 ; n4608
g4353 and n4607 n4608_not ; n4609
g4354 and n4515_not n4608_not ; n4610
g4355 and n4609_not n4610_not ; n4611
g4356 and n4350_not n4357_not ; n4612
g4357 and n4611 n4612 ; n4613
g4358 and n4611_not n4612_not ; n4614
g4359 and n4613_not n4614_not ; n4615
g4360 and b[20] n1302 ; n4616
g4361 and b[18] n1391 ; n4617
g4362 and b[19] n1297 ; n4618
g4363 and n4617_not n4618_not ; n4619
g4364 and n4616_not n4619 ; n4620
g4365 and n1305 n1846 ; n4621
g4366 and n4620 n4621_not ; n4622
g4367 and a[17] n4622_not ; n4623
g4368 and a[17] n4623_not ; n4624
g4369 and n4622_not n4623_not ; n4625
g4370 and n4624_not n4625_not ; n4626
g4371 and n4615 n4626_not ; n4627
g4372 and n4615_not n4626 ; n4628
g4373 and n4504_not n4628_not ; n4629
g4374 and n4627_not n4629 ; n4630
g4375 and n4504_not n4630_not ; n4631
g4376 and n4627_not n4630_not ; n4632
g4377 and n4628_not n4632 ; n4633
g4378 and n4631_not n4633_not ; n4634
g4379 and b[23] n951 ; n4635
g4380 and b[21] n1056 ; n4636
g4381 and b[22] n946 ; n4637
g4382 and n4636_not n4637_not ; n4638
g4383 and n4635_not n4638 ; n4639
g4384 and n954 n2300 ; n4640
g4385 and n4639 n4640_not ; n4641
g4386 and a[14] n4641_not ; n4642
g4387 and a[14] n4642_not ; n4643
g4388 and n4641_not n4642_not ; n4644
g4389 and n4643_not n4644_not ; n4645
g4390 and n4634 n4645 ; n4646
g4391 and n4634_not n4645_not ; n4647
g4392 and n4646_not n4647_not ; n4648
g4393 and n4503_not n4648 ; n4649
g4394 and n4503 n4648_not ; n4650
g4395 and n4649_not n4650_not ; n4651
g4396 and n4502 n4651_not ; n4652
g4397 and n4502_not n4651 ; n4653
g4398 and n4652_not n4653_not ; n4654
g4399 and n4414_not n4654 ; n4655
g4400 and n4414 n4654_not ; n4656
g4401 and n4655_not n4656_not ; n4657
g4402 and n4491_not n4657 ; n4658
g4403 and n4657 n4658_not ; n4659
g4404 and n4491_not n4658_not ; n4660
g4405 and n4659_not n4660_not ; n4661
g4406 and n4428_not n4434_not ; n4662
g4407 and n4661 n4662 ; n4663
g4408 and n4661_not n4662_not ; n4664
g4409 and n4663_not n4664_not ; n4665
g4410 and b[32] n362 ; n4666
g4411 and b[30] n403 ; n4667
g4412 and b[31] n357 ; n4668
g4413 and n4667_not n4668_not ; n4669
g4414 and n4666_not n4669 ; n4670
g4415 and n365 n4013 ; n4671
g4416 and n4670 n4671_not ; n4672
g4417 and a[5] n4672_not ; n4673
g4418 and a[5] n4673_not ; n4674
g4419 and n4672_not n4673_not ; n4675
g4420 and n4674_not n4675_not ; n4676
g4421 and n4665 n4676_not ; n4677
g4422 and n4665_not n4676 ; n4678
g4423 and n4452_not n4678_not ; n4679
g4424 and n4677_not n4679 ; n4680
g4425 and n4452_not n4680_not ; n4681
g4426 and n4677_not n4680_not ; n4682
g4427 and n4678_not n4682 ; n4683
g4428 and n4681_not n4683_not ; n4684
g4429 and b[35] n266 ; n4685
g4430 and b[33] n284 ; n4686
g4431 and b[34] n261 ; n4687
g4432 and n4686_not n4687_not ; n4688
g4433 and n4685_not n4688 ; n4689
g4434 and n4462_not n4464_not ; n4690
g4435 and b[34]_not b[35]_not ; n4691
g4436 and b[34] b[35] ; n4692
g4437 and n4691_not n4692_not ; n4693
g4438 and n4690_not n4693 ; n4694
g4439 and n4690 n4693_not ; n4695
g4440 and n4694_not n4695_not ; n4696
g4441 and n269 n4696 ; n4697
g4442 and n4689 n4697_not ; n4698
g4443 and a[2] n4698_not ; n4699
g4444 and a[2] n4699_not ; n4700
g4445 and n4698_not n4699_not ; n4701
g4446 and n4700_not n4701_not ; n4702
g4447 and n4684_not n4702 ; n4703
g4448 and n4684 n4702_not ; n4704
g4449 and n4703_not n4704_not ; n4705
g4450 and n4480_not n4705_not ; n4706
g4451 and n4480 n4705 ; n4707
g4452 and n4706_not n4707_not ; f[35]
g4453 and b[33] n362 ; n4709
g4454 and b[31] n403 ; n4710
g4455 and b[32] n357 ; n4711
g4456 and n4710_not n4711_not ; n4712
g4457 and n4709_not n4712 ; n4713
g4458 and n365 n4223 ; n4714
g4459 and n4713 n4714_not ; n4715
g4460 and a[5] n4715_not ; n4716
g4461 and a[5] n4716_not ; n4717
g4462 and n4715_not n4716_not ; n4718
g4463 and n4717_not n4718_not ; n4719
g4464 and n4658_not n4664_not ; n4720
g4465 and n4653_not n4655_not ; n4721
g4466 and b[27] n700 ; n4722
g4467 and b[25] n767 ; n4723
g4468 and b[26] n695 ; n4724
g4469 and n4723_not n4724_not ; n4725
g4470 and n4722_not n4725 ; n4726
g4471 and n703 n2990 ; n4727
g4472 and n4726 n4727_not ; n4728
g4473 and a[11] n4728_not ; n4729
g4474 and a[11] n4729_not ; n4730
g4475 and n4728_not n4729_not ; n4731
g4476 and n4730_not n4731_not ; n4732
g4477 and n4647_not n4649_not ; n4733
g4478 and n4608_not n4614_not ; n4734
g4479 and n4603_not n4605_not ; n4735
g4480 and b[15] n2048 ; n4736
g4481 and b[13] n2198 ; n4737
g4482 and b[14] n2043 ; n4738
g4483 and n4737_not n4738_not ; n4739
g4484 and n4736_not n4739 ; n4740
g4485 and n1131 n2051 ; n4741
g4486 and n4740 n4741_not ; n4742
g4487 and a[23] n4742_not ; n4743
g4488 and a[23] n4743_not ; n4744
g4489 and n4742_not n4743_not ; n4745
g4490 and n4744_not n4745_not ; n4746
g4491 and n4576_not n4580_not ; n4747
g4492 and b[6] n3638 ; n4748
g4493 and b[4] n3843 ; n4749
g4494 and b[5] n3633 ; n4750
g4495 and n4749_not n4750_not ; n4751
g4496 and n4748_not n4751 ; n4752
g4497 and n459 n3641 ; n4753
g4498 and n4752 n4753_not ; n4754
g4499 and a[32] n4754_not ; n4755
g4500 and a[32] n4755_not ; n4756
g4501 and n4754_not n4755_not ; n4757
g4502 and n4756_not n4757_not ; n4758
g4503 and a[35] a[36]_not ; n4759
g4504 and a[35]_not a[36] ; n4760
g4505 and n4759_not n4760_not ; n4761
g4506 and b[0] n4761_not ; n4762
g4507 and n4544_not n4762 ; n4763
g4508 and n4544 n4762_not ; n4764
g4509 and n4763_not n4764_not ; n4765
g4510 and b[3] n4287 ; n4766
g4511 and b[1] n4532 ; n4767
g4512 and b[2] n4282 ; n4768
g4513 and n4767_not n4768_not ; n4769
g4514 and n4766_not n4769 ; n4770
g4515 and n318 n4290 ; n4771
g4516 and n4770 n4771_not ; n4772
g4517 and a[35] n4772_not ; n4773
g4518 and a[35] n4773_not ; n4774
g4519 and n4772_not n4773_not ; n4775
g4520 and n4774_not n4775_not ; n4776
g4521 and n4765_not n4776_not ; n4777
g4522 and n4765 n4776 ; n4778
g4523 and n4777_not n4778_not ; n4779
g4524 and n4758_not n4779 ; n4780
g4525 and n4779 n4780_not ; n4781
g4526 and n4758_not n4780_not ; n4782
g4527 and n4781_not n4782_not ; n4783
g4528 and n4562_not n4783 ; n4784
g4529 and n4562 n4783_not ; n4785
g4530 and n4784_not n4785_not ; n4786
g4531 and b[9] n3050 ; n4787
g4532 and b[7] n3243 ; n4788
g4533 and b[8] n3045 ; n4789
g4534 and n4788_not n4789_not ; n4790
g4535 and n4787_not n4790 ; n4791
g4536 and n651 n3053 ; n4792
g4537 and n4791 n4792_not ; n4793
g4538 and a[29] n4793_not ; n4794
g4539 and a[29] n4794_not ; n4795
g4540 and n4793_not n4794_not ; n4796
g4541 and n4795_not n4796_not ; n4797
g4542 and n4786_not n4797_not ; n4798
g4543 and n4786 n4797 ; n4799
g4544 and n4798_not n4799_not ; n4800
g4545 and n4747 n4800_not ; n4801
g4546 and n4747_not n4800 ; n4802
g4547 and n4801_not n4802_not ; n4803
g4548 and b[12] n2539 ; n4804
g4549 and b[10] n2685 ; n4805
g4550 and b[11] n2534 ; n4806
g4551 and n4805_not n4806_not ; n4807
g4552 and n4804_not n4807 ; n4808
g4553 and n842 n2542 ; n4809
g4554 and n4808 n4809_not ; n4810
g4555 and a[26] n4810_not ; n4811
g4556 and a[26] n4811_not ; n4812
g4557 and n4810_not n4811_not ; n4813
g4558 and n4812_not n4813_not ; n4814
g4559 and n4803_not n4814 ; n4815
g4560 and n4803 n4814_not ; n4816
g4561 and n4815_not n4816_not ; n4817
g4562 and n4583_not n4587_not ; n4818
g4563 and n4817 n4818_not ; n4819
g4564 and n4817_not n4818 ; n4820
g4565 and n4819_not n4820_not ; n4821
g4566 and n4746_not n4821 ; n4822
g4567 and n4821 n4822_not ; n4823
g4568 and n4746_not n4822_not ; n4824
g4569 and n4823_not n4824_not ; n4825
g4570 and n4735_not n4825 ; n4826
g4571 and n4735 n4825_not ; n4827
g4572 and n4826_not n4827_not ; n4828
g4573 and b[18] n1627 ; n4829
g4574 and b[16] n1763 ; n4830
g4575 and b[17] n1622 ; n4831
g4576 and n4830_not n4831_not ; n4832
g4577 and n4829_not n4832 ; n4833
g4578 and n1566 n1630 ; n4834
g4579 and n4833 n4834_not ; n4835
g4580 and a[20] n4835_not ; n4836
g4581 and a[20] n4836_not ; n4837
g4582 and n4835_not n4836_not ; n4838
g4583 and n4837_not n4838_not ; n4839
g4584 and n4828_not n4839_not ; n4840
g4585 and n4828 n4839 ; n4841
g4586 and n4840_not n4841_not ; n4842
g4587 and n4734 n4842_not ; n4843
g4588 and n4734_not n4842 ; n4844
g4589 and n4843_not n4844_not ; n4845
g4590 and b[21] n1302 ; n4846
g4591 and b[19] n1391 ; n4847
g4592 and b[20] n1297 ; n4848
g4593 and n4847_not n4848_not ; n4849
g4594 and n4846_not n4849 ; n4850
g4595 and n1305 n1984 ; n4851
g4596 and n4850 n4851_not ; n4852
g4597 and a[17] n4852_not ; n4853
g4598 and a[17] n4853_not ; n4854
g4599 and n4852_not n4853_not ; n4855
g4600 and n4854_not n4855_not ; n4856
g4601 and n4845 n4856_not ; n4857
g4602 and n4845 n4857_not ; n4858
g4603 and n4856_not n4857_not ; n4859
g4604 and n4858_not n4859_not ; n4860
g4605 and n4632_not n4860 ; n4861
g4606 and n4632 n4860_not ; n4862
g4607 and n4861_not n4862_not ; n4863
g4608 and b[24] n951 ; n4864
g4609 and b[22] n1056 ; n4865
g4610 and b[23] n946 ; n4866
g4611 and n4865_not n4866_not ; n4867
g4612 and n4864_not n4867 ; n4868
g4613 and n954 n2458 ; n4869
g4614 and n4868 n4869_not ; n4870
g4615 and a[14] n4870_not ; n4871
g4616 and a[14] n4871_not ; n4872
g4617 and n4870_not n4871_not ; n4873
g4618 and n4872_not n4873_not ; n4874
g4619 and n4863 n4874 ; n4875
g4620 and n4863_not n4874_not ; n4876
g4621 and n4875_not n4876_not ; n4877
g4622 and n4733_not n4877 ; n4878
g4623 and n4733 n4877_not ; n4879
g4624 and n4878_not n4879_not ; n4880
g4625 and n4732_not n4880 ; n4881
g4626 and n4880 n4881_not ; n4882
g4627 and n4732_not n4881_not ; n4883
g4628 and n4882_not n4883_not ; n4884
g4629 and n4721_not n4884 ; n4885
g4630 and n4721 n4884_not ; n4886
g4631 and n4885_not n4886_not ; n4887
g4632 and b[30] n511 ; n4888
g4633 and b[28] n541 ; n4889
g4634 and b[29] n506 ; n4890
g4635 and n4889_not n4890_not ; n4891
g4636 and n4888_not n4891 ; n4892
g4637 and n514 n3577 ; n4893
g4638 and n4892 n4893_not ; n4894
g4639 and a[8] n4894_not ; n4895
g4640 and a[8] n4895_not ; n4896
g4641 and n4894_not n4895_not ; n4897
g4642 and n4896_not n4897_not ; n4898
g4643 and n4887 n4898 ; n4899
g4644 and n4887_not n4898_not ; n4900
g4645 and n4899_not n4900_not ; n4901
g4646 and n4720_not n4901 ; n4902
g4647 and n4720 n4901_not ; n4903
g4648 and n4902_not n4903_not ; n4904
g4649 and n4719_not n4904 ; n4905
g4650 and n4719 n4904_not ; n4906
g4651 and n4905_not n4906_not ; n4907
g4652 and n4682_not n4907 ; n4908
g4653 and n4682 n4907_not ; n4909
g4654 and n4908_not n4909_not ; n4910
g4655 and b[36] n266 ; n4911
g4656 and b[34] n284 ; n4912
g4657 and b[35] n261 ; n4913
g4658 and n4912_not n4913_not ; n4914
g4659 and n4911_not n4914 ; n4915
g4660 and n4692_not n4694_not ; n4916
g4661 and b[35]_not b[36]_not ; n4917
g4662 and b[35] b[36] ; n4918
g4663 and n4917_not n4918_not ; n4919
g4664 and n4916_not n4919 ; n4920
g4665 and n4916 n4919_not ; n4921
g4666 and n4920_not n4921_not ; n4922
g4667 and n269 n4922 ; n4923
g4668 and n4915 n4923_not ; n4924
g4669 and a[2] n4924_not ; n4925
g4670 and a[2] n4925_not ; n4926
g4671 and n4924_not n4925_not ; n4927
g4672 and n4926_not n4927_not ; n4928
g4673 and n4910 n4928_not ; n4929
g4674 and n4910 n4929_not ; n4930
g4675 and n4928_not n4929_not ; n4931
g4676 and n4930_not n4931_not ; n4932
g4677 and n4684_not n4702_not ; n4933
g4678 and n4706_not n4933_not ; n4934
g4679 and n4932_not n4934_not ; n4935
g4680 and n4932 n4934 ; n4936
g4681 and n4935_not n4936_not ; f[36]
g4682 and n4929_not n4935_not ; n4938
g4683 and b[34] n362 ; n4939
g4684 and b[32] n403 ; n4940
g4685 and b[33] n357 ; n4941
g4686 and n4940_not n4941_not ; n4942
g4687 and n4939_not n4942 ; n4943
g4688 and n365 n4466 ; n4944
g4689 and n4943 n4944_not ; n4945
g4690 and a[5] n4945_not ; n4946
g4691 and a[5] n4946_not ; n4947
g4692 and n4945_not n4946_not ; n4948
g4693 and n4947_not n4948_not ; n4949
g4694 and n4900_not n4902_not ; n4950
g4695 and b[31] n511 ; n4951
g4696 and b[29] n541 ; n4952
g4697 and b[30] n506 ; n4953
g4698 and n4952_not n4953_not ; n4954
g4699 and n4951_not n4954 ; n4955
g4700 and n514 n3796 ; n4956
g4701 and n4955 n4956_not ; n4957
g4702 and a[8] n4957_not ; n4958
g4703 and a[8] n4958_not ; n4959
g4704 and n4957_not n4958_not ; n4960
g4705 and n4959_not n4960_not ; n4961
g4706 and n4721_not n4884_not ; n4962
g4707 and n4881_not n4962_not ; n4963
g4708 and n4876_not n4878_not ; n4964
g4709 and b[16] n2048 ; n4965
g4710 and b[14] n2198 ; n4966
g4711 and b[15] n2043 ; n4967
g4712 and n4966_not n4967_not ; n4968
g4713 and n4965_not n4968 ; n4969
g4714 and n1237 n2051 ; n4970
g4715 and n4969 n4970_not ; n4971
g4716 and a[23] n4971_not ; n4972
g4717 and a[23] n4972_not ; n4973
g4718 and n4971_not n4972_not ; n4974
g4719 and n4973_not n4974_not ; n4975
g4720 and n4816_not n4819_not ; n4976
g4721 and b[13] n2539 ; n4977
g4722 and b[11] n2685 ; n4978
g4723 and b[12] n2534 ; n4979
g4724 and n4978_not n4979_not ; n4980
g4725 and n4977_not n4980 ; n4981
g4726 and n1008 n2542 ; n4982
g4727 and n4981 n4982_not ; n4983
g4728 and a[26] n4983_not ; n4984
g4729 and a[26] n4984_not ; n4985
g4730 and n4983_not n4984_not ; n4986
g4731 and n4985_not n4986_not ; n4987
g4732 and n4798_not n4802_not ; n4988
g4733 and b[10] n3050 ; n4989
g4734 and b[8] n3243 ; n4990
g4735 and b[9] n3045 ; n4991
g4736 and n4990_not n4991_not ; n4992
g4737 and n4989_not n4992 ; n4993
g4738 and n738 n3053 ; n4994
g4739 and n4993 n4994_not ; n4995
g4740 and a[29] n4995_not ; n4996
g4741 and a[29] n4996_not ; n4997
g4742 and n4995_not n4996_not ; n4998
g4743 and n4997_not n4998_not ; n4999
g4744 and n4562_not n4783_not ; n5000
g4745 and n4780_not n5000_not ; n5001
g4746 and b[7] n3638 ; n5002
g4747 and b[5] n3843 ; n5003
g4748 and b[6] n3633 ; n5004
g4749 and n5003_not n5004_not ; n5005
g4750 and n5002_not n5005 ; n5006
g4751 and n484 n3641 ; n5007
g4752 and n5006 n5007_not ; n5008
g4753 and a[32] n5008_not ; n5009
g4754 and a[32] n5009_not ; n5010
g4755 and n5008_not n5009_not ; n5011
g4756 and n5010_not n5011_not ; n5012
g4757 and n4544 n4762 ; n5013
g4758 and n4777_not n5013_not ; n5014
g4759 and b[4] n4287 ; n5015
g4760 and b[2] n4532 ; n5016
g4761 and b[3] n4282 ; n5017
g4762 and n5016_not n5017_not ; n5018
g4763 and n5015_not n5018 ; n5019
g4764 and n346 n4290 ; n5020
g4765 and n5019 n5020_not ; n5021
g4766 and a[35] n5021_not ; n5022
g4767 and a[35] n5022_not ; n5023
g4768 and n5021_not n5022_not ; n5024
g4769 and n5023_not n5024_not ; n5025
g4770 and a[38] n4762_not ; n5026
g4771 and a[36]_not a[37] ; n5027
g4772 and a[36] a[37]_not ; n5028
g4773 and n5027_not n5028_not ; n5029
g4774 and n4761 n5029_not ; n5030
g4775 and b[0] n5030 ; n5031
g4776 and a[37]_not a[38] ; n5032
g4777 and a[37] a[38]_not ; n5033
g4778 and n5032_not n5033_not ; n5034
g4779 and n4761_not n5034 ; n5035
g4780 and b[1] n5035 ; n5036
g4781 and n5031_not n5036_not ; n5037
g4782 and n4761_not n5034_not ; n5038
g4783 and n272_not n5038 ; n5039
g4784 and n5037 n5039_not ; n5040
g4785 and a[38] n5040_not ; n5041
g4786 and a[38] n5041_not ; n5042
g4787 and n5040_not n5041_not ; n5043
g4788 and n5042_not n5043_not ; n5044
g4789 and n5026 n5044_not ; n5045
g4790 and n5026_not n5044 ; n5046
g4791 and n5045_not n5046_not ; n5047
g4792 and n5025 n5047_not ; n5048
g4793 and n5025_not n5047 ; n5049
g4794 and n5048_not n5049_not ; n5050
g4795 and n5014_not n5050 ; n5051
g4796 and n5014 n5050_not ; n5052
g4797 and n5051_not n5052_not ; n5053
g4798 and n5012 n5053_not ; n5054
g4799 and n5012_not n5053 ; n5055
g4800 and n5054_not n5055_not ; n5056
g4801 and n5001_not n5056 ; n5057
g4802 and n5001 n5056_not ; n5058
g4803 and n5057_not n5058_not ; n5059
g4804 and n4999 n5059_not ; n5060
g4805 and n4999_not n5059 ; n5061
g4806 and n5060_not n5061_not ; n5062
g4807 and n4988_not n5062 ; n5063
g4808 and n4988 n5062_not ; n5064
g4809 and n5063_not n5064_not ; n5065
g4810 and n4987 n5065_not ; n5066
g4811 and n4987_not n5065 ; n5067
g4812 and n5066_not n5067_not ; n5068
g4813 and n4976_not n5068 ; n5069
g4814 and n4976 n5068_not ; n5070
g4815 and n5069_not n5070_not ; n5071
g4816 and n4975_not n5071 ; n5072
g4817 and n5071 n5072_not ; n5073
g4818 and n4975_not n5072_not ; n5074
g4819 and n5073_not n5074_not ; n5075
g4820 and n4735_not n4825_not ; n5076
g4821 and n4822_not n5076_not ; n5077
g4822 and n5075 n5077 ; n5078
g4823 and n5075_not n5077_not ; n5079
g4824 and n5078_not n5079_not ; n5080
g4825 and b[19] n1627 ; n5081
g4826 and b[17] n1763 ; n5082
g4827 and b[18] n1622 ; n5083
g4828 and n5082_not n5083_not ; n5084
g4829 and n5081_not n5084 ; n5085
g4830 and n1630 n1708 ; n5086
g4831 and n5085 n5086_not ; n5087
g4832 and a[20] n5087_not ; n5088
g4833 and a[20] n5088_not ; n5089
g4834 and n5087_not n5088_not ; n5090
g4835 and n5089_not n5090_not ; n5091
g4836 and n5080 n5091_not ; n5092
g4837 and n5080 n5092_not ; n5093
g4838 and n5091_not n5092_not ; n5094
g4839 and n5093_not n5094_not ; n5095
g4840 and n4840_not n4844_not ; n5096
g4841 and n5095 n5096 ; n5097
g4842 and n5095_not n5096_not ; n5098
g4843 and n5097_not n5098_not ; n5099
g4844 and b[22] n1302 ; n5100
g4845 and b[20] n1391 ; n5101
g4846 and b[21] n1297 ; n5102
g4847 and n5101_not n5102_not ; n5103
g4848 and n5100_not n5103 ; n5104
g4849 and n1305 n2145 ; n5105
g4850 and n5104 n5105_not ; n5106
g4851 and a[17] n5106_not ; n5107
g4852 and a[17] n5107_not ; n5108
g4853 and n5106_not n5107_not ; n5109
g4854 and n5108_not n5109_not ; n5110
g4855 and n5099 n5110_not ; n5111
g4856 and n5099 n5111_not ; n5112
g4857 and n5110_not n5111_not ; n5113
g4858 and n5112_not n5113_not ; n5114
g4859 and n4632_not n4860_not ; n5115
g4860 and n4857_not n5115_not ; n5116
g4861 and n5114 n5116 ; n5117
g4862 and n5114_not n5116_not ; n5118
g4863 and n5117_not n5118_not ; n5119
g4864 and b[25] n951 ; n5120
g4865 and b[23] n1056 ; n5121
g4866 and b[24] n946 ; n5122
g4867 and n5121_not n5122_not ; n5123
g4868 and n5120_not n5123 ; n5124
g4869 and n954 n2485 ; n5125
g4870 and n5124 n5125_not ; n5126
g4871 and a[14] n5126_not ; n5127
g4872 and a[14] n5127_not ; n5128
g4873 and n5126_not n5127_not ; n5129
g4874 and n5128_not n5129_not ; n5130
g4875 and n5119 n5130_not ; n5131
g4876 and n5119_not n5130 ; n5132
g4877 and n4964_not n5132_not ; n5133
g4878 and n5131_not n5133 ; n5134
g4879 and n4964_not n5134_not ; n5135
g4880 and n5131_not n5134_not ; n5136
g4881 and n5132_not n5136 ; n5137
g4882 and n5135_not n5137_not ; n5138
g4883 and b[28] n700 ; n5139
g4884 and b[26] n767 ; n5140
g4885 and b[27] n695 ; n5141
g4886 and n5140_not n5141_not ; n5142
g4887 and n5139_not n5142 ; n5143
g4888 and n703 n3189 ; n5144
g4889 and n5143 n5144_not ; n5145
g4890 and a[11] n5145_not ; n5146
g4891 and a[11] n5146_not ; n5147
g4892 and n5145_not n5146_not ; n5148
g4893 and n5147_not n5148_not ; n5149
g4894 and n5138 n5149 ; n5150
g4895 and n5138_not n5149_not ; n5151
g4896 and n5150_not n5151_not ; n5152
g4897 and n4963_not n5152 ; n5153
g4898 and n4963 n5152_not ; n5154
g4899 and n5153_not n5154_not ; n5155
g4900 and n4961 n5155_not ; n5156
g4901 and n4961_not n5155 ; n5157
g4902 and n5156_not n5157_not ; n5158
g4903 and n4950_not n5158 ; n5159
g4904 and n4950 n5158_not ; n5160
g4905 and n5159_not n5160_not ; n5161
g4906 and n4949_not n5161 ; n5162
g4907 and n5161 n5162_not ; n5163
g4908 and n4949_not n5162_not ; n5164
g4909 and n5163_not n5164_not ; n5165
g4910 and n4905_not n4908_not ; n5166
g4911 and n5165 n5166 ; n5167
g4912 and n5165_not n5166_not ; n5168
g4913 and n5167_not n5168_not ; n5169
g4914 and b[37] n266 ; n5170
g4915 and b[35] n284 ; n5171
g4916 and b[36] n261 ; n5172
g4917 and n5171_not n5172_not ; n5173
g4918 and n5170_not n5173 ; n5174
g4919 and n4918_not n4920_not ; n5175
g4920 and b[36]_not b[37]_not ; n5176
g4921 and b[36] b[37] ; n5177
g4922 and n5176_not n5177_not ; n5178
g4923 and n5175_not n5178 ; n5179
g4924 and n5175 n5178_not ; n5180
g4925 and n5179_not n5180_not ; n5181
g4926 and n269 n5181 ; n5182
g4927 and n5174 n5182_not ; n5183
g4928 and a[2] n5183_not ; n5184
g4929 and a[2] n5184_not ; n5185
g4930 and n5183_not n5184_not ; n5186
g4931 and n5185_not n5186_not ; n5187
g4932 and n5169_not n5187 ; n5188
g4933 and n5169 n5187_not ; n5189
g4934 and n5188_not n5189_not ; n5190
g4935 and n4938_not n5190 ; n5191
g4936 and n4938 n5190_not ; n5192
g4937 and n5191_not n5192_not ; f[37]
g4938 and b[38] n266 ; n5194
g4939 and b[36] n284 ; n5195
g4940 and b[37] n261 ; n5196
g4941 and n5195_not n5196_not ; n5197
g4942 and n5194_not n5197 ; n5198
g4943 and n5177_not n5179_not ; n5199
g4944 and b[37]_not b[38]_not ; n5200
g4945 and b[37] b[38] ; n5201
g4946 and n5200_not n5201_not ; n5202
g4947 and n5199_not n5202 ; n5203
g4948 and n5199 n5202_not ; n5204
g4949 and n5203_not n5204_not ; n5205
g4950 and n269 n5205 ; n5206
g4951 and n5198 n5206_not ; n5207
g4952 and a[2] n5207_not ; n5208
g4953 and a[2] n5208_not ; n5209
g4954 and n5207_not n5208_not ; n5210
g4955 and n5209_not n5210_not ; n5211
g4956 and n5162_not n5168_not ; n5212
g4957 and b[35] n362 ; n5213
g4958 and b[33] n403 ; n5214
g4959 and b[34] n357 ; n5215
g4960 and n5214_not n5215_not ; n5216
g4961 and n5213_not n5216 ; n5217
g4962 and n365 n4696 ; n5218
g4963 and n5217 n5218_not ; n5219
g4964 and a[5] n5219_not ; n5220
g4965 and a[5] n5220_not ; n5221
g4966 and n5219_not n5220_not ; n5222
g4967 and n5221_not n5222_not ; n5223
g4968 and n5157_not n5159_not ; n5224
g4969 and b[32] n511 ; n5225
g4970 and b[30] n541 ; n5226
g4971 and b[31] n506 ; n5227
g4972 and n5226_not n5227_not ; n5228
g4973 and n5225_not n5228 ; n5229
g4974 and n514 n4013 ; n5230
g4975 and n5229 n5230_not ; n5231
g4976 and a[8] n5231_not ; n5232
g4977 and a[8] n5232_not ; n5233
g4978 and n5231_not n5232_not ; n5234
g4979 and n5233_not n5234_not ; n5235
g4980 and n5151_not n5153_not ; n5236
g4981 and b[29] n700 ; n5237
g4982 and b[27] n767 ; n5238
g4983 and b[28] n695 ; n5239
g4984 and n5238_not n5239_not ; n5240
g4985 and n5237_not n5240 ; n5241
g4986 and n703 n3383 ; n5242
g4987 and n5241 n5242_not ; n5243
g4988 and a[11] n5243_not ; n5244
g4989 and a[11] n5244_not ; n5245
g4990 and n5243_not n5244_not ; n5246
g4991 and n5245_not n5246_not ; n5247
g4992 and n5111_not n5118_not ; n5248
g4993 and b[17] n2048 ; n5249
g4994 and b[15] n2198 ; n5250
g4995 and b[16] n2043 ; n5251
g4996 and n5250_not n5251_not ; n5252
g4997 and n5249_not n5252 ; n5253
g4998 and n1356 n2051 ; n5254
g4999 and n5253 n5254_not ; n5255
g5000 and a[23] n5255_not ; n5256
g5001 and a[23] n5256_not ; n5257
g5002 and n5255_not n5256_not ; n5258
g5003 and n5257_not n5258_not ; n5259
g5004 and n5067_not n5069_not ; n5260
g5005 and n5061_not n5063_not ; n5261
g5006 and b[11] n3050 ; n5262
g5007 and b[9] n3243 ; n5263
g5008 and b[10] n3045 ; n5264
g5009 and n5263_not n5264_not ; n5265
g5010 and n5262_not n5265 ; n5266
g5011 and n818 n3053 ; n5267
g5012 and n5266 n5267_not ; n5268
g5013 and a[29] n5268_not ; n5269
g5014 and a[29] n5269_not ; n5270
g5015 and n5268_not n5269_not ; n5271
g5016 and n5270_not n5271_not ; n5272
g5017 and n5055_not n5057_not ; n5273
g5018 and n5049_not n5051_not ; n5274
g5019 and b[2] n5035 ; n5275
g5020 and n4761 n5034_not ; n5276
g5021 and n5029 n5276 ; n5277
g5022 and b[0] n5277 ; n5278
g5023 and b[1] n5030 ; n5279
g5024 and n5278_not n5279_not ; n5280
g5025 and n5275_not n5280 ; n5281
g5026 and n296 n5038 ; n5282
g5027 and n5281 n5282_not ; n5283
g5028 and a[38] n5283_not ; n5284
g5029 and a[38] n5284_not ; n5285
g5030 and n5283_not n5284_not ; n5286
g5031 and n5285_not n5286_not ; n5287
g5032 and n5045_not n5287 ; n5288
g5033 and n5045 n5287_not ; n5289
g5034 and n5288_not n5289_not ; n5290
g5035 and b[5] n4287 ; n5291
g5036 and b[3] n4532 ; n5292
g5037 and b[4] n4282 ; n5293
g5038 and n5292_not n5293_not ; n5294
g5039 and n5291_not n5294 ; n5295
g5040 and n394 n4290 ; n5296
g5041 and n5295 n5296_not ; n5297
g5042 and a[35] n5297_not ; n5298
g5043 and a[35] n5298_not ; n5299
g5044 and n5297_not n5298_not ; n5300
g5045 and n5299_not n5300_not ; n5301
g5046 and n5290 n5301_not ; n5302
g5047 and n5290 n5302_not ; n5303
g5048 and n5301_not n5302_not ; n5304
g5049 and n5303_not n5304_not ; n5305
g5050 and n5274_not n5305 ; n5306
g5051 and n5274 n5305_not ; n5307
g5052 and n5306_not n5307_not ; n5308
g5053 and b[8] n3638 ; n5309
g5054 and b[6] n3843 ; n5310
g5055 and b[7] n3633 ; n5311
g5056 and n5310_not n5311_not ; n5312
g5057 and n5309_not n5312 ; n5313
g5058 and n585 n3641 ; n5314
g5059 and n5313 n5314_not ; n5315
g5060 and a[32] n5315_not ; n5316
g5061 and a[32] n5316_not ; n5317
g5062 and n5315_not n5316_not ; n5318
g5063 and n5317_not n5318_not ; n5319
g5064 and n5308_not n5319_not ; n5320
g5065 and n5308 n5319 ; n5321
g5066 and n5320_not n5321_not ; n5322
g5067 and n5273_not n5322 ; n5323
g5068 and n5273 n5322_not ; n5324
g5069 and n5323_not n5324_not ; n5325
g5070 and n5272_not n5325 ; n5326
g5071 and n5272_not n5326_not ; n5327
g5072 and n5325 n5326_not ; n5328
g5073 and n5327_not n5328_not ; n5329
g5074 and n5261_not n5329_not ; n5330
g5075 and n5261_not n5330_not ; n5331
g5076 and n5329_not n5330_not ; n5332
g5077 and n5331_not n5332_not ; n5333
g5078 and b[14] n2539 ; n5334
g5079 and b[12] n2685 ; n5335
g5080 and b[13] n2534 ; n5336
g5081 and n5335_not n5336_not ; n5337
g5082 and n5334_not n5337 ; n5338
g5083 and n1034 n2542 ; n5339
g5084 and n5338 n5339_not ; n5340
g5085 and a[26] n5340_not ; n5341
g5086 and a[26] n5341_not ; n5342
g5087 and n5340_not n5341_not ; n5343
g5088 and n5342_not n5343_not ; n5344
g5089 and n5333 n5344 ; n5345
g5090 and n5333_not n5344_not ; n5346
g5091 and n5345_not n5346_not ; n5347
g5092 and n5260_not n5347 ; n5348
g5093 and n5260 n5347_not ; n5349
g5094 and n5348_not n5349_not ; n5350
g5095 and n5259_not n5350 ; n5351
g5096 and n5350 n5351_not ; n5352
g5097 and n5259_not n5351_not ; n5353
g5098 and n5352_not n5353_not ; n5354
g5099 and n5072_not n5079_not ; n5355
g5100 and n5354 n5355 ; n5356
g5101 and n5354_not n5355_not ; n5357
g5102 and n5356_not n5357_not ; n5358
g5103 and b[20] n1627 ; n5359
g5104 and b[18] n1763 ; n5360
g5105 and b[19] n1622 ; n5361
g5106 and n5360_not n5361_not ; n5362
g5107 and n5359_not n5362 ; n5363
g5108 and n1630 n1846 ; n5364
g5109 and n5363 n5364_not ; n5365
g5110 and a[20] n5365_not ; n5366
g5111 and a[20] n5366_not ; n5367
g5112 and n5365_not n5366_not ; n5368
g5113 and n5367_not n5368_not ; n5369
g5114 and n5358 n5369_not ; n5370
g5115 and n5358 n5370_not ; n5371
g5116 and n5369_not n5370_not ; n5372
g5117 and n5371_not n5372_not ; n5373
g5118 and n5092_not n5098_not ; n5374
g5119 and n5373 n5374 ; n5375
g5120 and n5373_not n5374_not ; n5376
g5121 and n5375_not n5376_not ; n5377
g5122 and b[23] n1302 ; n5378
g5123 and b[21] n1391 ; n5379
g5124 and b[22] n1297 ; n5380
g5125 and n5379_not n5380_not ; n5381
g5126 and n5378_not n5381 ; n5382
g5127 and n1305 n2300 ; n5383
g5128 and n5382 n5383_not ; n5384
g5129 and a[17] n5384_not ; n5385
g5130 and a[17] n5385_not ; n5386
g5131 and n5384_not n5385_not ; n5387
g5132 and n5386_not n5387_not ; n5388
g5133 and n5377 n5388_not ; n5389
g5134 and n5377_not n5388 ; n5390
g5135 and n5248_not n5390_not ; n5391
g5136 and n5389_not n5391 ; n5392
g5137 and n5248_not n5392_not ; n5393
g5138 and n5389_not n5392_not ; n5394
g5139 and n5390_not n5394 ; n5395
g5140 and n5393_not n5395_not ; n5396
g5141 and b[26] n951 ; n5397
g5142 and b[24] n1056 ; n5398
g5143 and b[25] n946 ; n5399
g5144 and n5398_not n5399_not ; n5400
g5145 and n5397_not n5400 ; n5401
g5146 and n954 n2813 ; n5402
g5147 and n5401 n5402_not ; n5403
g5148 and a[14] n5403_not ; n5404
g5149 and a[14] n5404_not ; n5405
g5150 and n5403_not n5404_not ; n5406
g5151 and n5405_not n5406_not ; n5407
g5152 and n5396 n5407 ; n5408
g5153 and n5396_not n5407_not ; n5409
g5154 and n5408_not n5409_not ; n5410
g5155 and n5136_not n5410 ; n5411
g5156 and n5136 n5410_not ; n5412
g5157 and n5411_not n5412_not ; n5413
g5158 and n5247 n5413_not ; n5414
g5159 and n5247_not n5413 ; n5415
g5160 and n5414_not n5415_not ; n5416
g5161 and n5236_not n5416 ; n5417
g5162 and n5236 n5416_not ; n5418
g5163 and n5417_not n5418_not ; n5419
g5164 and n5235 n5419_not ; n5420
g5165 and n5235_not n5419 ; n5421
g5166 and n5420_not n5421_not ; n5422
g5167 and n5224_not n5422 ; n5423
g5168 and n5224 n5422_not ; n5424
g5169 and n5423_not n5424_not ; n5425
g5170 and n5223 n5425_not ; n5426
g5171 and n5223_not n5425 ; n5427
g5172 and n5426_not n5427_not ; n5428
g5173 and n5212_not n5428 ; n5429
g5174 and n5212 n5428_not ; n5430
g5175 and n5429_not n5430_not ; n5431
g5176 and n5211_not n5431 ; n5432
g5177 and n5431 n5432_not ; n5433
g5178 and n5211_not n5432_not ; n5434
g5179 and n5433_not n5434_not ; n5435
g5180 and n5189_not n5191_not ; n5436
g5181 and n5435_not n5436_not ; n5437
g5182 and n5435 n5436 ; n5438
g5183 and n5437_not n5438_not ; f[38]
g5184 and b[39] n266 ; n5440
g5185 and b[37] n284 ; n5441
g5186 and b[38] n261 ; n5442
g5187 and n5441_not n5442_not ; n5443
g5188 and n5440_not n5443 ; n5444
g5189 and n5201_not n5203_not ; n5445
g5190 and b[38]_not b[39]_not ; n5446
g5191 and b[38] b[39] ; n5447
g5192 and n5446_not n5447_not ; n5448
g5193 and n5445_not n5448 ; n5449
g5194 and n5445 n5448_not ; n5450
g5195 and n5449_not n5450_not ; n5451
g5196 and n269 n5451 ; n5452
g5197 and n5444 n5452_not ; n5453
g5198 and a[2] n5453_not ; n5454
g5199 and a[2] n5454_not ; n5455
g5200 and n5453_not n5454_not ; n5456
g5201 and n5455_not n5456_not ; n5457
g5202 and n5427_not n5429_not ; n5458
g5203 and n5421_not n5423_not ; n5459
g5204 and b[33] n511 ; n5460
g5205 and b[31] n541 ; n5461
g5206 and b[32] n506 ; n5462
g5207 and n5461_not n5462_not ; n5463
g5208 and n5460_not n5463 ; n5464
g5209 and n514 n4223 ; n5465
g5210 and n5464 n5465_not ; n5466
g5211 and a[8] n5466_not ; n5467
g5212 and a[8] n5467_not ; n5468
g5213 and n5466_not n5467_not ; n5469
g5214 and n5468_not n5469_not ; n5470
g5215 and n5415_not n5417_not ; n5471
g5216 and n5409_not n5411_not ; n5472
g5217 and b[27] n951 ; n5473
g5218 and b[25] n1056 ; n5474
g5219 and b[26] n946 ; n5475
g5220 and n5474_not n5475_not ; n5476
g5221 and n5473_not n5476 ; n5477
g5222 and n954 n2990 ; n5478
g5223 and n5477 n5478_not ; n5479
g5224 and a[14] n5479_not ; n5480
g5225 and a[14] n5480_not ; n5481
g5226 and n5479_not n5480_not ; n5482
g5227 and n5481_not n5482_not ; n5483
g5228 and n5351_not n5357_not ; n5484
g5229 and n5346_not n5348_not ; n5485
g5230 and b[15] n2539 ; n5486
g5231 and b[13] n2685 ; n5487
g5232 and b[14] n2534 ; n5488
g5233 and n5487_not n5488_not ; n5489
g5234 and n5486_not n5489 ; n5490
g5235 and n1131 n2542 ; n5491
g5236 and n5490 n5491_not ; n5492
g5237 and a[26] n5492_not ; n5493
g5238 and a[26] n5493_not ; n5494
g5239 and n5492_not n5493_not ; n5495
g5240 and n5494_not n5495_not ; n5496
g5241 and b[6] n4287 ; n5497
g5242 and b[4] n4532 ; n5498
g5243 and b[5] n4282 ; n5499
g5244 and n5498_not n5499_not ; n5500
g5245 and n5497_not n5500 ; n5501
g5246 and n459 n4290 ; n5502
g5247 and n5501 n5502_not ; n5503
g5248 and a[35] n5503_not ; n5504
g5249 and a[35] n5504_not ; n5505
g5250 and n5503_not n5504_not ; n5506
g5251 and n5505_not n5506_not ; n5507
g5252 and a[38] a[39]_not ; n5508
g5253 and a[38]_not a[39] ; n5509
g5254 and n5508_not n5509_not ; n5510
g5255 and b[0] n5510_not ; n5511
g5256 and n5289_not n5511 ; n5512
g5257 and n5289 n5511_not ; n5513
g5258 and n5512_not n5513_not ; n5514
g5259 and b[3] n5035 ; n5515
g5260 and b[1] n5277 ; n5516
g5261 and b[2] n5030 ; n5517
g5262 and n5516_not n5517_not ; n5518
g5263 and n5515_not n5518 ; n5519
g5264 and n318 n5038 ; n5520
g5265 and n5519 n5520_not ; n5521
g5266 and a[38] n5521_not ; n5522
g5267 and a[38] n5522_not ; n5523
g5268 and n5521_not n5522_not ; n5524
g5269 and n5523_not n5524_not ; n5525
g5270 and n5514_not n5525_not ; n5526
g5271 and n5514 n5525 ; n5527
g5272 and n5526_not n5527_not ; n5528
g5273 and n5507_not n5528 ; n5529
g5274 and n5528 n5529_not ; n5530
g5275 and n5507_not n5529_not ; n5531
g5276 and n5530_not n5531_not ; n5532
g5277 and n5274_not n5305_not ; n5533
g5278 and n5302_not n5533_not ; n5534
g5279 and n5532 n5534 ; n5535
g5280 and n5532_not n5534_not ; n5536
g5281 and n5535_not n5536_not ; n5537
g5282 and b[9] n3638 ; n5538
g5283 and b[7] n3843 ; n5539
g5284 and b[8] n3633 ; n5540
g5285 and n5539_not n5540_not ; n5541
g5286 and n5538_not n5541 ; n5542
g5287 and n651 n3641 ; n5543
g5288 and n5542 n5543_not ; n5544
g5289 and a[32] n5544_not ; n5545
g5290 and a[32] n5545_not ; n5546
g5291 and n5544_not n5545_not ; n5547
g5292 and n5546_not n5547_not ; n5548
g5293 and n5537 n5548_not ; n5549
g5294 and n5537 n5549_not ; n5550
g5295 and n5548_not n5549_not ; n5551
g5296 and n5550_not n5551_not ; n5552
g5297 and n5320_not n5323_not ; n5553
g5298 and n5552 n5553 ; n5554
g5299 and n5552_not n5553_not ; n5555
g5300 and n5554_not n5555_not ; n5556
g5301 and b[12] n3050 ; n5557
g5302 and b[10] n3243 ; n5558
g5303 and b[11] n3045 ; n5559
g5304 and n5558_not n5559_not ; n5560
g5305 and n5557_not n5560 ; n5561
g5306 and n842 n3053 ; n5562
g5307 and n5561 n5562_not ; n5563
g5308 and a[29] n5563_not ; n5564
g5309 and a[29] n5564_not ; n5565
g5310 and n5563_not n5564_not ; n5566
g5311 and n5565_not n5566_not ; n5567
g5312 and n5556_not n5567 ; n5568
g5313 and n5556 n5567_not ; n5569
g5314 and n5568_not n5569_not ; n5570
g5315 and n5326_not n5330_not ; n5571
g5316 and n5570 n5571_not ; n5572
g5317 and n5570_not n5571 ; n5573
g5318 and n5572_not n5573_not ; n5574
g5319 and n5496_not n5574 ; n5575
g5320 and n5574 n5575_not ; n5576
g5321 and n5496_not n5575_not ; n5577
g5322 and n5576_not n5577_not ; n5578
g5323 and n5485_not n5578 ; n5579
g5324 and n5485 n5578_not ; n5580
g5325 and n5579_not n5580_not ; n5581
g5326 and b[18] n2048 ; n5582
g5327 and b[16] n2198 ; n5583
g5328 and b[17] n2043 ; n5584
g5329 and n5583_not n5584_not ; n5585
g5330 and n5582_not n5585 ; n5586
g5331 and n1566 n2051 ; n5587
g5332 and n5586 n5587_not ; n5588
g5333 and a[23] n5588_not ; n5589
g5334 and a[23] n5589_not ; n5590
g5335 and n5588_not n5589_not ; n5591
g5336 and n5590_not n5591_not ; n5592
g5337 and n5581_not n5592_not ; n5593
g5338 and n5581 n5592 ; n5594
g5339 and n5593_not n5594_not ; n5595
g5340 and n5484 n5595_not ; n5596
g5341 and n5484_not n5595 ; n5597
g5342 and n5596_not n5597_not ; n5598
g5343 and b[21] n1627 ; n5599
g5344 and b[19] n1763 ; n5600
g5345 and b[20] n1622 ; n5601
g5346 and n5600_not n5601_not ; n5602
g5347 and n5599_not n5602 ; n5603
g5348 and n1630 n1984 ; n5604
g5349 and n5603 n5604_not ; n5605
g5350 and a[20] n5605_not ; n5606
g5351 and a[20] n5606_not ; n5607
g5352 and n5605_not n5606_not ; n5608
g5353 and n5607_not n5608_not ; n5609
g5354 and n5598 n5609_not ; n5610
g5355 and n5598 n5610_not ; n5611
g5356 and n5609_not n5610_not ; n5612
g5357 and n5611_not n5612_not ; n5613
g5358 and n5370_not n5376_not ; n5614
g5359 and n5613 n5614 ; n5615
g5360 and n5613_not n5614_not ; n5616
g5361 and n5615_not n5616_not ; n5617
g5362 and b[24] n1302 ; n5618
g5363 and b[22] n1391 ; n5619
g5364 and b[23] n1297 ; n5620
g5365 and n5619_not n5620_not ; n5621
g5366 and n5618_not n5621 ; n5622
g5367 and n1305 n2458 ; n5623
g5368 and n5622 n5623_not ; n5624
g5369 and a[17] n5624_not ; n5625
g5370 and a[17] n5625_not ; n5626
g5371 and n5624_not n5625_not ; n5627
g5372 and n5626_not n5627_not ; n5628
g5373 and n5617_not n5628 ; n5629
g5374 and n5617 n5628_not ; n5630
g5375 and n5629_not n5630_not ; n5631
g5376 and n5394_not n5631 ; n5632
g5377 and n5394 n5631_not ; n5633
g5378 and n5632_not n5633_not ; n5634
g5379 and n5483_not n5634 ; n5635
g5380 and n5634 n5635_not ; n5636
g5381 and n5483_not n5635_not ; n5637
g5382 and n5636_not n5637_not ; n5638
g5383 and n5472_not n5638 ; n5639
g5384 and n5472 n5638_not ; n5640
g5385 and n5639_not n5640_not ; n5641
g5386 and b[30] n700 ; n5642
g5387 and b[28] n767 ; n5643
g5388 and b[29] n695 ; n5644
g5389 and n5643_not n5644_not ; n5645
g5390 and n5642_not n5645 ; n5646
g5391 and n703 n3577 ; n5647
g5392 and n5646 n5647_not ; n5648
g5393 and a[11] n5648_not ; n5649
g5394 and a[11] n5649_not ; n5650
g5395 and n5648_not n5649_not ; n5651
g5396 and n5650_not n5651_not ; n5652
g5397 and n5641_not n5652_not ; n5653
g5398 and n5641 n5652 ; n5654
g5399 and n5653_not n5654_not ; n5655
g5400 and n5471_not n5655 ; n5656
g5401 and n5471 n5655_not ; n5657
g5402 and n5656_not n5657_not ; n5658
g5403 and n5470_not n5658 ; n5659
g5404 and n5658 n5659_not ; n5660
g5405 and n5470_not n5659_not ; n5661
g5406 and n5660_not n5661_not ; n5662
g5407 and n5459_not n5662 ; n5663
g5408 and n5459 n5662_not ; n5664
g5409 and n5663_not n5664_not ; n5665
g5410 and b[36] n362 ; n5666
g5411 and b[34] n403 ; n5667
g5412 and b[35] n357 ; n5668
g5413 and n5667_not n5668_not ; n5669
g5414 and n5666_not n5669 ; n5670
g5415 and n365 n4922 ; n5671
g5416 and n5670 n5671_not ; n5672
g5417 and a[5] n5672_not ; n5673
g5418 and a[5] n5673_not ; n5674
g5419 and n5672_not n5673_not ; n5675
g5420 and n5674_not n5675_not ; n5676
g5421 and n5665 n5676 ; n5677
g5422 and n5665_not n5676_not ; n5678
g5423 and n5677_not n5678_not ; n5679
g5424 and n5458_not n5679 ; n5680
g5425 and n5458 n5679_not ; n5681
g5426 and n5680_not n5681_not ; n5682
g5427 and n5457_not n5682 ; n5683
g5428 and n5682 n5683_not ; n5684
g5429 and n5457_not n5683_not ; n5685
g5430 and n5684_not n5685_not ; n5686
g5431 and n5432_not n5437_not ; n5687
g5432 and n5686_not n5687_not ; n5688
g5433 and n5686 n5687 ; n5689
g5434 and n5688_not n5689_not ; f[39]
g5435 and n5683_not n5688_not ; n5691
g5436 and n5678_not n5680_not ; n5692
g5437 and b[37] n362 ; n5693
g5438 and b[35] n403 ; n5694
g5439 and b[36] n357 ; n5695
g5440 and n5694_not n5695_not ; n5696
g5441 and n5693_not n5696 ; n5697
g5442 and n365 n5181 ; n5698
g5443 and n5697 n5698_not ; n5699
g5444 and a[5] n5699_not ; n5700
g5445 and a[5] n5700_not ; n5701
g5446 and n5699_not n5700_not ; n5702
g5447 and n5701_not n5702_not ; n5703
g5448 and n5459_not n5662_not ; n5704
g5449 and n5659_not n5704_not ; n5705
g5450 and b[34] n511 ; n5706
g5451 and b[32] n541 ; n5707
g5452 and b[33] n506 ; n5708
g5453 and n5707_not n5708_not ; n5709
g5454 and n5706_not n5709 ; n5710
g5455 and n514 n4466 ; n5711
g5456 and n5710 n5711_not ; n5712
g5457 and a[8] n5712_not ; n5713
g5458 and a[8] n5713_not ; n5714
g5459 and n5712_not n5713_not ; n5715
g5460 and n5714_not n5715_not ; n5716
g5461 and n5653_not n5656_not ; n5717
g5462 and n5472_not n5638_not ; n5718
g5463 and n5635_not n5718_not ; n5719
g5464 and b[28] n951 ; n5720
g5465 and b[26] n1056 ; n5721
g5466 and b[27] n946 ; n5722
g5467 and n5721_not n5722_not ; n5723
g5468 and n5720_not n5723 ; n5724
g5469 and n954 n3189 ; n5725
g5470 and n5724 n5725_not ; n5726
g5471 and a[14] n5726_not ; n5727
g5472 and a[14] n5727_not ; n5728
g5473 and n5726_not n5727_not ; n5729
g5474 and n5728_not n5729_not ; n5730
g5475 and b[16] n2539 ; n5731
g5476 and b[14] n2685 ; n5732
g5477 and b[15] n2534 ; n5733
g5478 and n5732_not n5733_not ; n5734
g5479 and n5731_not n5734 ; n5735
g5480 and n1237 n2542 ; n5736
g5481 and n5735 n5736_not ; n5737
g5482 and a[26] n5737_not ; n5738
g5483 and a[26] n5738_not ; n5739
g5484 and n5737_not n5738_not ; n5740
g5485 and n5739_not n5740_not ; n5741
g5486 and n5569_not n5572_not ; n5742
g5487 and n5549_not n5555_not ; n5743
g5488 and b[7] n4287 ; n5744
g5489 and b[5] n4532 ; n5745
g5490 and b[6] n4282 ; n5746
g5491 and n5745_not n5746_not ; n5747
g5492 and n5744_not n5747 ; n5748
g5493 and n484 n4290 ; n5749
g5494 and n5748 n5749_not ; n5750
g5495 and a[35] n5750_not ; n5751
g5496 and a[35] n5751_not ; n5752
g5497 and n5750_not n5751_not ; n5753
g5498 and n5752_not n5753_not ; n5754
g5499 and n5289 n5511 ; n5755
g5500 and n5526_not n5755_not ; n5756
g5501 and b[4] n5035 ; n5757
g5502 and b[2] n5277 ; n5758
g5503 and b[3] n5030 ; n5759
g5504 and n5758_not n5759_not ; n5760
g5505 and n5757_not n5760 ; n5761
g5506 and n346 n5038 ; n5762
g5507 and n5761 n5762_not ; n5763
g5508 and a[38] n5763_not ; n5764
g5509 and a[38] n5764_not ; n5765
g5510 and n5763_not n5764_not ; n5766
g5511 and n5765_not n5766_not ; n5767
g5512 and a[41] n5511_not ; n5768
g5513 and a[39]_not a[40] ; n5769
g5514 and a[39] a[40]_not ; n5770
g5515 and n5769_not n5770_not ; n5771
g5516 and n5510 n5771_not ; n5772
g5517 and b[0] n5772 ; n5773
g5518 and a[40]_not a[41] ; n5774
g5519 and a[40] a[41]_not ; n5775
g5520 and n5774_not n5775_not ; n5776
g5521 and n5510_not n5776 ; n5777
g5522 and b[1] n5777 ; n5778
g5523 and n5773_not n5778_not ; n5779
g5524 and n5510_not n5776_not ; n5780
g5525 and n272_not n5780 ; n5781
g5526 and n5779 n5781_not ; n5782
g5527 and a[41] n5782_not ; n5783
g5528 and a[41] n5783_not ; n5784
g5529 and n5782_not n5783_not ; n5785
g5530 and n5784_not n5785_not ; n5786
g5531 and n5768 n5786_not ; n5787
g5532 and n5768_not n5786 ; n5788
g5533 and n5787_not n5788_not ; n5789
g5534 and n5767 n5789_not ; n5790
g5535 and n5767_not n5789 ; n5791
g5536 and n5790_not n5791_not ; n5792
g5537 and n5756_not n5792 ; n5793
g5538 and n5756 n5792_not ; n5794
g5539 and n5793_not n5794_not ; n5795
g5540 and n5754_not n5795 ; n5796
g5541 and n5795 n5796_not ; n5797
g5542 and n5754_not n5796_not ; n5798
g5543 and n5797_not n5798_not ; n5799
g5544 and n5529_not n5536_not ; n5800
g5545 and n5799 n5800 ; n5801
g5546 and n5799_not n5800_not ; n5802
g5547 and n5801_not n5802_not ; n5803
g5548 and b[10] n3638 ; n5804
g5549 and b[8] n3843 ; n5805
g5550 and b[9] n3633 ; n5806
g5551 and n5805_not n5806_not ; n5807
g5552 and n5804_not n5807 ; n5808
g5553 and n738 n3641 ; n5809
g5554 and n5808 n5809_not ; n5810
g5555 and a[32] n5810_not ; n5811
g5556 and a[32] n5811_not ; n5812
g5557 and n5810_not n5811_not ; n5813
g5558 and n5812_not n5813_not ; n5814
g5559 and n5803 n5814_not ; n5815
g5560 and n5803_not n5814 ; n5816
g5561 and n5743_not n5816_not ; n5817
g5562 and n5815_not n5817 ; n5818
g5563 and n5743_not n5818_not ; n5819
g5564 and n5815_not n5818_not ; n5820
g5565 and n5816_not n5820 ; n5821
g5566 and n5819_not n5821_not ; n5822
g5567 and b[13] n3050 ; n5823
g5568 and b[11] n3243 ; n5824
g5569 and b[12] n3045 ; n5825
g5570 and n5824_not n5825_not ; n5826
g5571 and n5823_not n5826 ; n5827
g5572 and n1008 n3053 ; n5828
g5573 and n5827 n5828_not ; n5829
g5574 and a[29] n5829_not ; n5830
g5575 and a[29] n5830_not ; n5831
g5576 and n5829_not n5830_not ; n5832
g5577 and n5831_not n5832_not ; n5833
g5578 and n5822 n5833 ; n5834
g5579 and n5822_not n5833_not ; n5835
g5580 and n5834_not n5835_not ; n5836
g5581 and n5742_not n5836 ; n5837
g5582 and n5742 n5836_not ; n5838
g5583 and n5837_not n5838_not ; n5839
g5584 and n5741_not n5839 ; n5840
g5585 and n5839 n5840_not ; n5841
g5586 and n5741_not n5840_not ; n5842
g5587 and n5841_not n5842_not ; n5843
g5588 and n5485_not n5578_not ; n5844
g5589 and n5575_not n5844_not ; n5845
g5590 and n5843 n5845 ; n5846
g5591 and n5843_not n5845_not ; n5847
g5592 and n5846_not n5847_not ; n5848
g5593 and b[19] n2048 ; n5849
g5594 and b[17] n2198 ; n5850
g5595 and b[18] n2043 ; n5851
g5596 and n5850_not n5851_not ; n5852
g5597 and n5849_not n5852 ; n5853
g5598 and n1708 n2051 ; n5854
g5599 and n5853 n5854_not ; n5855
g5600 and a[23] n5855_not ; n5856
g5601 and a[23] n5856_not ; n5857
g5602 and n5855_not n5856_not ; n5858
g5603 and n5857_not n5858_not ; n5859
g5604 and n5848 n5859_not ; n5860
g5605 and n5848 n5860_not ; n5861
g5606 and n5859_not n5860_not ; n5862
g5607 and n5861_not n5862_not ; n5863
g5608 and n5593_not n5597_not ; n5864
g5609 and n5863 n5864 ; n5865
g5610 and n5863_not n5864_not ; n5866
g5611 and n5865_not n5866_not ; n5867
g5612 and b[22] n1627 ; n5868
g5613 and b[20] n1763 ; n5869
g5614 and b[21] n1622 ; n5870
g5615 and n5869_not n5870_not ; n5871
g5616 and n5868_not n5871 ; n5872
g5617 and n1630 n2145 ; n5873
g5618 and n5872 n5873_not ; n5874
g5619 and a[20] n5874_not ; n5875
g5620 and a[20] n5875_not ; n5876
g5621 and n5874_not n5875_not ; n5877
g5622 and n5876_not n5877_not ; n5878
g5623 and n5867 n5878_not ; n5879
g5624 and n5867 n5879_not ; n5880
g5625 and n5878_not n5879_not ; n5881
g5626 and n5880_not n5881_not ; n5882
g5627 and n5610_not n5616_not ; n5883
g5628 and n5882 n5883 ; n5884
g5629 and n5882_not n5883_not ; n5885
g5630 and n5884_not n5885_not ; n5886
g5631 and b[25] n1302 ; n5887
g5632 and b[23] n1391 ; n5888
g5633 and b[24] n1297 ; n5889
g5634 and n5888_not n5889_not ; n5890
g5635 and n5887_not n5890 ; n5891
g5636 and n1305 n2485 ; n5892
g5637 and n5891 n5892_not ; n5893
g5638 and a[17] n5893_not ; n5894
g5639 and a[17] n5894_not ; n5895
g5640 and n5893_not n5894_not ; n5896
g5641 and n5895_not n5896_not ; n5897
g5642 and n5886 n5897_not ; n5898
g5643 and n5886 n5898_not ; n5899
g5644 and n5897_not n5898_not ; n5900
g5645 and n5899_not n5900_not ; n5901
g5646 and n5630_not n5632_not ; n5902
g5647 and n5901_not n5902_not ; n5903
g5648 and n5901 n5902 ; n5904
g5649 and n5903_not n5904_not ; n5905
g5650 and n5730_not n5905 ; n5906
g5651 and n5730_not n5906_not ; n5907
g5652 and n5905 n5906_not ; n5908
g5653 and n5907_not n5908_not ; n5909
g5654 and n5719_not n5909_not ; n5910
g5655 and n5719_not n5910_not ; n5911
g5656 and n5909_not n5910_not ; n5912
g5657 and n5911_not n5912_not ; n5913
g5658 and b[31] n700 ; n5914
g5659 and b[29] n767 ; n5915
g5660 and b[30] n695 ; n5916
g5661 and n5915_not n5916_not ; n5917
g5662 and n5914_not n5917 ; n5918
g5663 and n703 n3796 ; n5919
g5664 and n5918 n5919_not ; n5920
g5665 and a[11] n5920_not ; n5921
g5666 and a[11] n5921_not ; n5922
g5667 and n5920_not n5921_not ; n5923
g5668 and n5922_not n5923_not ; n5924
g5669 and n5913 n5924 ; n5925
g5670 and n5913_not n5924_not ; n5926
g5671 and n5925_not n5926_not ; n5927
g5672 and n5717_not n5927 ; n5928
g5673 and n5717 n5927_not ; n5929
g5674 and n5928_not n5929_not ; n5930
g5675 and n5716 n5930_not ; n5931
g5676 and n5716_not n5930 ; n5932
g5677 and n5931_not n5932_not ; n5933
g5678 and n5705_not n5933 ; n5934
g5679 and n5705 n5933_not ; n5935
g5680 and n5934_not n5935_not ; n5936
g5681 and n5703_not n5936 ; n5937
g5682 and n5936 n5937_not ; n5938
g5683 and n5703_not n5937_not ; n5939
g5684 and n5938_not n5939_not ; n5940
g5685 and n5692_not n5940 ; n5941
g5686 and n5692 n5940_not ; n5942
g5687 and n5941_not n5942_not ; n5943
g5688 and b[40] n266 ; n5944
g5689 and b[38] n284 ; n5945
g5690 and b[39] n261 ; n5946
g5691 and n5945_not n5946_not ; n5947
g5692 and n5944_not n5947 ; n5948
g5693 and n5447_not n5449_not ; n5949
g5694 and b[39]_not b[40]_not ; n5950
g5695 and b[39] b[40] ; n5951
g5696 and n5950_not n5951_not ; n5952
g5697 and n5949_not n5952 ; n5953
g5698 and n5949 n5952_not ; n5954
g5699 and n5953_not n5954_not ; n5955
g5700 and n269 n5955 ; n5956
g5701 and n5948 n5956_not ; n5957
g5702 and a[2] n5957_not ; n5958
g5703 and a[2] n5958_not ; n5959
g5704 and n5957_not n5958_not ; n5960
g5705 and n5959_not n5960_not ; n5961
g5706 and n5943_not n5961_not ; n5962
g5707 and n5943 n5961 ; n5963
g5708 and n5962_not n5963_not ; n5964
g5709 and n5691_not n5964 ; n5965
g5710 and n5691 n5964_not ; n5966
g5711 and n5965_not n5966_not ; f[40]
g5712 and n5962_not n5965_not ; n5968
g5713 and n5692_not n5940_not ; n5969
g5714 and n5937_not n5969_not ; n5970
g5715 and n5932_not n5934_not ; n5971
g5716 and b[35] n511 ; n5972
g5717 and b[33] n541 ; n5973
g5718 and b[34] n506 ; n5974
g5719 and n5973_not n5974_not ; n5975
g5720 and n5972_not n5975 ; n5976
g5721 and n514 n4696 ; n5977
g5722 and n5976 n5977_not ; n5978
g5723 and a[8] n5978_not ; n5979
g5724 and a[8] n5979_not ; n5980
g5725 and n5978_not n5979_not ; n5981
g5726 and n5980_not n5981_not ; n5982
g5727 and n5926_not n5928_not ; n5983
g5728 and b[32] n700 ; n5984
g5729 and b[30] n767 ; n5985
g5730 and b[31] n695 ; n5986
g5731 and n5985_not n5986_not ; n5987
g5732 and n5984_not n5987 ; n5988
g5733 and n703 n4013 ; n5989
g5734 and n5988 n5989_not ; n5990
g5735 and a[11] n5990_not ; n5991
g5736 and a[11] n5991_not ; n5992
g5737 and n5990_not n5991_not ; n5993
g5738 and n5992_not n5993_not ; n5994
g5739 and n5906_not n5910_not ; n5995
g5740 and b[29] n951 ; n5996
g5741 and b[27] n1056 ; n5997
g5742 and b[28] n946 ; n5998
g5743 and n5997_not n5998_not ; n5999
g5744 and n5996_not n5999 ; n6000
g5745 and n954 n3383 ; n6001
g5746 and n6000 n6001_not ; n6002
g5747 and a[14] n6002_not ; n6003
g5748 and a[14] n6003_not ; n6004
g5749 and n6002_not n6003_not ; n6005
g5750 and n6004_not n6005_not ; n6006
g5751 and n5898_not n5903_not ; n6007
g5752 and n5879_not n5885_not ; n6008
g5753 and b[20] n2048 ; n6009
g5754 and b[18] n2198 ; n6010
g5755 and b[19] n2043 ; n6011
g5756 and n6010_not n6011_not ; n6012
g5757 and n6009_not n6012 ; n6013
g5758 and n1846 n2051 ; n6014
g5759 and n6013 n6014_not ; n6015
g5760 and a[23] n6015_not ; n6016
g5761 and a[23] n6016_not ; n6017
g5762 and n6015_not n6016_not ; n6018
g5763 and n6017_not n6018_not ; n6019
g5764 and n5840_not n5847_not ; n6020
g5765 and b[17] n2539 ; n6021
g5766 and b[15] n2685 ; n6022
g5767 and b[16] n2534 ; n6023
g5768 and n6022_not n6023_not ; n6024
g5769 and n6021_not n6024 ; n6025
g5770 and n1356 n2542 ; n6026
g5771 and n6025 n6026_not ; n6027
g5772 and a[26] n6027_not ; n6028
g5773 and a[26] n6028_not ; n6029
g5774 and n6027_not n6028_not ; n6030
g5775 and n6029_not n6030_not ; n6031
g5776 and n5835_not n5837_not ; n6032
g5777 and b[14] n3050 ; n6033
g5778 and b[12] n3243 ; n6034
g5779 and b[13] n3045 ; n6035
g5780 and n6034_not n6035_not ; n6036
g5781 and n6033_not n6036 ; n6037
g5782 and n1034 n3053 ; n6038
g5783 and n6037 n6038_not ; n6039
g5784 and a[29] n6039_not ; n6040
g5785 and a[29] n6040_not ; n6041
g5786 and n6039_not n6040_not ; n6042
g5787 and n6041_not n6042_not ; n6043
g5788 and n5796_not n5802_not ; n6044
g5789 and b[8] n4287 ; n6045
g5790 and b[6] n4532 ; n6046
g5791 and b[7] n4282 ; n6047
g5792 and n6046_not n6047_not ; n6048
g5793 and n6045_not n6048 ; n6049
g5794 and n585 n4290 ; n6050
g5795 and n6049 n6050_not ; n6051
g5796 and a[35] n6051_not ; n6052
g5797 and a[35] n6052_not ; n6053
g5798 and n6051_not n6052_not ; n6054
g5799 and n6053_not n6054_not ; n6055
g5800 and n5791_not n5793_not ; n6056
g5801 and b[2] n5777 ; n6057
g5802 and n5510 n5776_not ; n6058
g5803 and n5771 n6058 ; n6059
g5804 and b[0] n6059 ; n6060
g5805 and b[1] n5772 ; n6061
g5806 and n6060_not n6061_not ; n6062
g5807 and n6057_not n6062 ; n6063
g5808 and n296 n5780 ; n6064
g5809 and n6063 n6064_not ; n6065
g5810 and a[41] n6065_not ; n6066
g5811 and a[41] n6066_not ; n6067
g5812 and n6065_not n6066_not ; n6068
g5813 and n6067_not n6068_not ; n6069
g5814 and n5787_not n6069 ; n6070
g5815 and n5787 n6069_not ; n6071
g5816 and n6070_not n6071_not ; n6072
g5817 and b[5] n5035 ; n6073
g5818 and b[3] n5277 ; n6074
g5819 and b[4] n5030 ; n6075
g5820 and n6074_not n6075_not ; n6076
g5821 and n6073_not n6076 ; n6077
g5822 and n394 n5038 ; n6078
g5823 and n6077 n6078_not ; n6079
g5824 and a[38] n6079_not ; n6080
g5825 and a[38] n6080_not ; n6081
g5826 and n6079_not n6080_not ; n6082
g5827 and n6081_not n6082_not ; n6083
g5828 and n6072 n6083_not ; n6084
g5829 and n6072 n6084_not ; n6085
g5830 and n6083_not n6084_not ; n6086
g5831 and n6085_not n6086_not ; n6087
g5832 and n6056_not n6087_not ; n6088
g5833 and n6056 n6087 ; n6089
g5834 and n6088_not n6089_not ; n6090
g5835 and n6055_not n6090 ; n6091
g5836 and n6055_not n6091_not ; n6092
g5837 and n6090 n6091_not ; n6093
g5838 and n6092_not n6093_not ; n6094
g5839 and n6044_not n6094_not ; n6095
g5840 and n6044_not n6095_not ; n6096
g5841 and n6094_not n6095_not ; n6097
g5842 and n6096_not n6097_not ; n6098
g5843 and b[11] n3638 ; n6099
g5844 and b[9] n3843 ; n6100
g5845 and b[10] n3633 ; n6101
g5846 and n6100_not n6101_not ; n6102
g5847 and n6099_not n6102 ; n6103
g5848 and n818 n3641 ; n6104
g5849 and n6103 n6104_not ; n6105
g5850 and a[32] n6105_not ; n6106
g5851 and a[32] n6106_not ; n6107
g5852 and n6105_not n6106_not ; n6108
g5853 and n6107_not n6108_not ; n6109
g5854 and n6098 n6109 ; n6110
g5855 and n6098_not n6109_not ; n6111
g5856 and n6110_not n6111_not ; n6112
g5857 and n5820_not n6112 ; n6113
g5858 and n5820 n6112_not ; n6114
g5859 and n6113_not n6114_not ; n6115
g5860 and n6043 n6115_not ; n6116
g5861 and n6043_not n6115 ; n6117
g5862 and n6116_not n6117_not ; n6118
g5863 and n6032_not n6118 ; n6119
g5864 and n6032 n6118_not ; n6120
g5865 and n6119_not n6120_not ; n6121
g5866 and n6031 n6121_not ; n6122
g5867 and n6031_not n6121 ; n6123
g5868 and n6122_not n6123_not ; n6124
g5869 and n6020_not n6124 ; n6125
g5870 and n6020 n6124_not ; n6126
g5871 and n6125_not n6126_not ; n6127
g5872 and n6019_not n6127 ; n6128
g5873 and n6127 n6128_not ; n6129
g5874 and n6019_not n6128_not ; n6130
g5875 and n6129_not n6130_not ; n6131
g5876 and n5860_not n5866_not ; n6132
g5877 and n6131 n6132 ; n6133
g5878 and n6131_not n6132_not ; n6134
g5879 and n6133_not n6134_not ; n6135
g5880 and b[23] n1627 ; n6136
g5881 and b[21] n1763 ; n6137
g5882 and b[22] n1622 ; n6138
g5883 and n6137_not n6138_not ; n6139
g5884 and n6136_not n6139 ; n6140
g5885 and n1630 n2300 ; n6141
g5886 and n6140 n6141_not ; n6142
g5887 and a[20] n6142_not ; n6143
g5888 and a[20] n6143_not ; n6144
g5889 and n6142_not n6143_not ; n6145
g5890 and n6144_not n6145_not ; n6146
g5891 and n6135 n6146_not ; n6147
g5892 and n6135_not n6146 ; n6148
g5893 and n6008_not n6148_not ; n6149
g5894 and n6147_not n6149 ; n6150
g5895 and n6008_not n6150_not ; n6151
g5896 and n6147_not n6150_not ; n6152
g5897 and n6148_not n6152 ; n6153
g5898 and n6151_not n6153_not ; n6154
g5899 and b[26] n1302 ; n6155
g5900 and b[24] n1391 ; n6156
g5901 and b[25] n1297 ; n6157
g5902 and n6156_not n6157_not ; n6158
g5903 and n6155_not n6158 ; n6159
g5904 and n1305 n2813 ; n6160
g5905 and n6159 n6160_not ; n6161
g5906 and a[17] n6161_not ; n6162
g5907 and a[17] n6162_not ; n6163
g5908 and n6161_not n6162_not ; n6164
g5909 and n6163_not n6164_not ; n6165
g5910 and n6154 n6165 ; n6166
g5911 and n6154_not n6165_not ; n6167
g5912 and n6166_not n6167_not ; n6168
g5913 and n6007_not n6168 ; n6169
g5914 and n6007 n6168_not ; n6170
g5915 and n6169_not n6170_not ; n6171
g5916 and n6006 n6171_not ; n6172
g5917 and n6006_not n6171 ; n6173
g5918 and n6172_not n6173_not ; n6174
g5919 and n5995_not n6174 ; n6175
g5920 and n5995 n6174_not ; n6176
g5921 and n6175_not n6176_not ; n6177
g5922 and n5994 n6177_not ; n6178
g5923 and n5994_not n6177 ; n6179
g5924 and n6178_not n6179_not ; n6180
g5925 and n5983_not n6180 ; n6181
g5926 and n5983 n6180_not ; n6182
g5927 and n6181_not n6182_not ; n6183
g5928 and n5982_not n6183 ; n6184
g5929 and n6183 n6184_not ; n6185
g5930 and n5982_not n6184_not ; n6186
g5931 and n6185_not n6186_not ; n6187
g5932 and n5971_not n6187 ; n6188
g5933 and n5971 n6187_not ; n6189
g5934 and n6188_not n6189_not ; n6190
g5935 and b[38] n362 ; n6191
g5936 and b[36] n403 ; n6192
g5937 and b[37] n357 ; n6193
g5938 and n6192_not n6193_not ; n6194
g5939 and n6191_not n6194 ; n6195
g5940 and n365 n5205 ; n6196
g5941 and n6195 n6196_not ; n6197
g5942 and a[5] n6197_not ; n6198
g5943 and a[5] n6198_not ; n6199
g5944 and n6197_not n6198_not ; n6200
g5945 and n6199_not n6200_not ; n6201
g5946 and n6190_not n6201_not ; n6202
g5947 and n6190 n6201 ; n6203
g5948 and n6202_not n6203_not ; n6204
g5949 and n5970 n6204_not ; n6205
g5950 and n5970_not n6204 ; n6206
g5951 and n6205_not n6206_not ; n6207
g5952 and b[41] n266 ; n6208
g5953 and b[39] n284 ; n6209
g5954 and b[40] n261 ; n6210
g5955 and n6209_not n6210_not ; n6211
g5956 and n6208_not n6211 ; n6212
g5957 and n5951_not n5953_not ; n6213
g5958 and b[40]_not b[41]_not ; n6214
g5959 and b[40] b[41] ; n6215
g5960 and n6214_not n6215_not ; n6216
g5961 and n6213_not n6216 ; n6217
g5962 and n6213 n6216_not ; n6218
g5963 and n6217_not n6218_not ; n6219
g5964 and n269 n6219 ; n6220
g5965 and n6212 n6220_not ; n6221
g5966 and a[2] n6221_not ; n6222
g5967 and a[2] n6222_not ; n6223
g5968 and n6221_not n6222_not ; n6224
g5969 and n6223_not n6224_not ; n6225
g5970 and n6207_not n6225 ; n6226
g5971 and n6207 n6225_not ; n6227
g5972 and n6226_not n6227_not ; n6228
g5973 and n5968_not n6228 ; n6229
g5974 and n5968 n6228_not ; n6230
g5975 and n6229_not n6230_not ; f[41]
g5976 and n6202_not n6206_not ; n6232
g5977 and b[39] n362 ; n6233
g5978 and b[37] n403 ; n6234
g5979 and b[38] n357 ; n6235
g5980 and n6234_not n6235_not ; n6236
g5981 and n6233_not n6236 ; n6237
g5982 and n365 n5451 ; n6238
g5983 and n6237 n6238_not ; n6239
g5984 and a[5] n6239_not ; n6240
g5985 and a[5] n6240_not ; n6241
g5986 and n6239_not n6240_not ; n6242
g5987 and n6241_not n6242_not ; n6243
g5988 and n5971_not n6187_not ; n6244
g5989 and n6184_not n6244_not ; n6245
g5990 and n6179_not n6181_not ; n6246
g5991 and b[33] n700 ; n6247
g5992 and b[31] n767 ; n6248
g5993 and b[32] n695 ; n6249
g5994 and n6248_not n6249_not ; n6250
g5995 and n6247_not n6250 ; n6251
g5996 and n703 n4223 ; n6252
g5997 and n6251 n6252_not ; n6253
g5998 and a[11] n6253_not ; n6254
g5999 and a[11] n6254_not ; n6255
g6000 and n6253_not n6254_not ; n6256
g6001 and n6255_not n6256_not ; n6257
g6002 and n6173_not n6175_not ; n6258
g6003 and n6167_not n6169_not ; n6259
g6004 and b[27] n1302 ; n6260
g6005 and b[25] n1391 ; n6261
g6006 and b[26] n1297 ; n6262
g6007 and n6261_not n6262_not ; n6263
g6008 and n6260_not n6263 ; n6264
g6009 and n1305 n2990 ; n6265
g6010 and n6264 n6265_not ; n6266
g6011 and a[17] n6266_not ; n6267
g6012 and a[17] n6267_not ; n6268
g6013 and n6266_not n6267_not ; n6269
g6014 and n6268_not n6269_not ; n6270
g6015 and b[21] n2048 ; n6271
g6016 and b[19] n2198 ; n6272
g6017 and b[20] n2043 ; n6273
g6018 and n6272_not n6273_not ; n6274
g6019 and n6271_not n6274 ; n6275
g6020 and n1984 n2051 ; n6276
g6021 and n6275 n6276_not ; n6277
g6022 and a[23] n6277_not ; n6278
g6023 and a[23] n6278_not ; n6279
g6024 and n6277_not n6278_not ; n6280
g6025 and n6279_not n6280_not ; n6281
g6026 and n6123_not n6125_not ; n6282
g6027 and n6117_not n6119_not ; n6283
g6028 and n6111_not n6113_not ; n6284
g6029 and b[12] n3638 ; n6285
g6030 and b[10] n3843 ; n6286
g6031 and b[11] n3633 ; n6287
g6032 and n6286_not n6287_not ; n6288
g6033 and n6285_not n6288 ; n6289
g6034 and n842 n3641 ; n6290
g6035 and n6289 n6290_not ; n6291
g6036 and a[32] n6291_not ; n6292
g6037 and a[32] n6292_not ; n6293
g6038 and n6291_not n6292_not ; n6294
g6039 and n6293_not n6294_not ; n6295
g6040 and n6091_not n6095_not ; n6296
g6041 and b[6] n5035 ; n6297
g6042 and b[4] n5277 ; n6298
g6043 and b[5] n5030 ; n6299
g6044 and n6298_not n6299_not ; n6300
g6045 and n6297_not n6300 ; n6301
g6046 and n459 n5038 ; n6302
g6047 and n6301 n6302_not ; n6303
g6048 and a[38] n6303_not ; n6304
g6049 and a[38] n6304_not ; n6305
g6050 and n6303_not n6304_not ; n6306
g6051 and n6305_not n6306_not ; n6307
g6052 and a[41] a[42]_not ; n6308
g6053 and a[41]_not a[42] ; n6309
g6054 and n6308_not n6309_not ; n6310
g6055 and b[0] n6310_not ; n6311
g6056 and n6071_not n6311 ; n6312
g6057 and n6071 n6311_not ; n6313
g6058 and n6312_not n6313_not ; n6314
g6059 and b[3] n5777 ; n6315
g6060 and b[1] n6059 ; n6316
g6061 and b[2] n5772 ; n6317
g6062 and n6316_not n6317_not ; n6318
g6063 and n6315_not n6318 ; n6319
g6064 and n318 n5780 ; n6320
g6065 and n6319 n6320_not ; n6321
g6066 and a[41] n6321_not ; n6322
g6067 and a[41] n6322_not ; n6323
g6068 and n6321_not n6322_not ; n6324
g6069 and n6323_not n6324_not ; n6325
g6070 and n6314_not n6325_not ; n6326
g6071 and n6314 n6325 ; n6327
g6072 and n6326_not n6327_not ; n6328
g6073 and n6307_not n6328 ; n6329
g6074 and n6328 n6329_not ; n6330
g6075 and n6307_not n6329_not ; n6331
g6076 and n6330_not n6331_not ; n6332
g6077 and n6084_not n6088_not ; n6333
g6078 and n6332 n6333 ; n6334
g6079 and n6332_not n6333_not ; n6335
g6080 and n6334_not n6335_not ; n6336
g6081 and b[9] n4287 ; n6337
g6082 and b[7] n4532 ; n6338
g6083 and b[8] n4282 ; n6339
g6084 and n6338_not n6339_not ; n6340
g6085 and n6337_not n6340 ; n6341
g6086 and n651 n4290 ; n6342
g6087 and n6341 n6342_not ; n6343
g6088 and a[35] n6343_not ; n6344
g6089 and a[35] n6344_not ; n6345
g6090 and n6343_not n6344_not ; n6346
g6091 and n6345_not n6346_not ; n6347
g6092 and n6336_not n6347 ; n6348
g6093 and n6336 n6347_not ; n6349
g6094 and n6348_not n6349_not ; n6350
g6095 and n6296_not n6350 ; n6351
g6096 and n6296 n6350_not ; n6352
g6097 and n6351_not n6352_not ; n6353
g6098 and n6295_not n6353 ; n6354
g6099 and n6295_not n6354_not ; n6355
g6100 and n6353 n6354_not ; n6356
g6101 and n6355_not n6356_not ; n6357
g6102 and n6284_not n6357_not ; n6358
g6103 and n6284_not n6358_not ; n6359
g6104 and n6357_not n6358_not ; n6360
g6105 and n6359_not n6360_not ; n6361
g6106 and b[15] n3050 ; n6362
g6107 and b[13] n3243 ; n6363
g6108 and b[14] n3045 ; n6364
g6109 and n6363_not n6364_not ; n6365
g6110 and n6362_not n6365 ; n6366
g6111 and n1131 n3053 ; n6367
g6112 and n6366 n6367_not ; n6368
g6113 and a[29] n6368_not ; n6369
g6114 and a[29] n6369_not ; n6370
g6115 and n6368_not n6369_not ; n6371
g6116 and n6370_not n6371_not ; n6372
g6117 and n6361_not n6372_not ; n6373
g6118 and n6361_not n6373_not ; n6374
g6119 and n6372_not n6373_not ; n6375
g6120 and n6374_not n6375_not ; n6376
g6121 and n6283_not n6376 ; n6377
g6122 and n6283 n6376_not ; n6378
g6123 and n6377_not n6378_not ; n6379
g6124 and b[18] n2539 ; n6380
g6125 and b[16] n2685 ; n6381
g6126 and b[17] n2534 ; n6382
g6127 and n6381_not n6382_not ; n6383
g6128 and n6380_not n6383 ; n6384
g6129 and n1566 n2542 ; n6385
g6130 and n6384 n6385_not ; n6386
g6131 and a[26] n6386_not ; n6387
g6132 and a[26] n6387_not ; n6388
g6133 and n6386_not n6387_not ; n6389
g6134 and n6388_not n6389_not ; n6390
g6135 and n6379_not n6390_not ; n6391
g6136 and n6379 n6390 ; n6392
g6137 and n6391_not n6392_not ; n6393
g6138 and n6282_not n6393 ; n6394
g6139 and n6282 n6393_not ; n6395
g6140 and n6394_not n6395_not ; n6396
g6141 and n6281_not n6396 ; n6397
g6142 and n6396 n6397_not ; n6398
g6143 and n6281_not n6397_not ; n6399
g6144 and n6398_not n6399_not ; n6400
g6145 and n6128_not n6134_not ; n6401
g6146 and n6400 n6401 ; n6402
g6147 and n6400_not n6401_not ; n6403
g6148 and n6402_not n6403_not ; n6404
g6149 and b[24] n1627 ; n6405
g6150 and b[22] n1763 ; n6406
g6151 and b[23] n1622 ; n6407
g6152 and n6406_not n6407_not ; n6408
g6153 and n6405_not n6408 ; n6409
g6154 and n1630 n2458 ; n6410
g6155 and n6409 n6410_not ; n6411
g6156 and a[20] n6411_not ; n6412
g6157 and a[20] n6412_not ; n6413
g6158 and n6411_not n6412_not ; n6414
g6159 and n6413_not n6414_not ; n6415
g6160 and n6404_not n6415 ; n6416
g6161 and n6404 n6415_not ; n6417
g6162 and n6416_not n6417_not ; n6418
g6163 and n6152_not n6418 ; n6419
g6164 and n6152 n6418_not ; n6420
g6165 and n6419_not n6420_not ; n6421
g6166 and n6270_not n6421 ; n6422
g6167 and n6421 n6422_not ; n6423
g6168 and n6270_not n6422_not ; n6424
g6169 and n6423_not n6424_not ; n6425
g6170 and n6259_not n6425 ; n6426
g6171 and n6259 n6425_not ; n6427
g6172 and n6426_not n6427_not ; n6428
g6173 and b[30] n951 ; n6429
g6174 and b[28] n1056 ; n6430
g6175 and b[29] n946 ; n6431
g6176 and n6430_not n6431_not ; n6432
g6177 and n6429_not n6432 ; n6433
g6178 and n954 n3577 ; n6434
g6179 and n6433 n6434_not ; n6435
g6180 and a[14] n6435_not ; n6436
g6181 and a[14] n6436_not ; n6437
g6182 and n6435_not n6436_not ; n6438
g6183 and n6437_not n6438_not ; n6439
g6184 and n6428_not n6439_not ; n6440
g6185 and n6428 n6439 ; n6441
g6186 and n6440_not n6441_not ; n6442
g6187 and n6258_not n6442 ; n6443
g6188 and n6258 n6442_not ; n6444
g6189 and n6443_not n6444_not ; n6445
g6190 and n6257_not n6445 ; n6446
g6191 and n6445 n6446_not ; n6447
g6192 and n6257_not n6446_not ; n6448
g6193 and n6447_not n6448_not ; n6449
g6194 and n6246_not n6449 ; n6450
g6195 and n6246 n6449_not ; n6451
g6196 and n6450_not n6451_not ; n6452
g6197 and b[36] n511 ; n6453
g6198 and b[34] n541 ; n6454
g6199 and b[35] n506 ; n6455
g6200 and n6454_not n6455_not ; n6456
g6201 and n6453_not n6456 ; n6457
g6202 and n514 n4922 ; n6458
g6203 and n6457 n6458_not ; n6459
g6204 and a[8] n6459_not ; n6460
g6205 and a[8] n6460_not ; n6461
g6206 and n6459_not n6460_not ; n6462
g6207 and n6461_not n6462_not ; n6463
g6208 and n6452 n6463 ; n6464
g6209 and n6452_not n6463_not ; n6465
g6210 and n6464_not n6465_not ; n6466
g6211 and n6245_not n6466 ; n6467
g6212 and n6245 n6466_not ; n6468
g6213 and n6467_not n6468_not ; n6469
g6214 and n6243_not n6469 ; n6470
g6215 and n6243_not n6470_not ; n6471
g6216 and n6469 n6470_not ; n6472
g6217 and n6471_not n6472_not ; n6473
g6218 and n6232_not n6473_not ; n6474
g6219 and n6232_not n6474_not ; n6475
g6220 and n6473_not n6474_not ; n6476
g6221 and n6475_not n6476_not ; n6477
g6222 and b[42] n266 ; n6478
g6223 and b[40] n284 ; n6479
g6224 and b[41] n261 ; n6480
g6225 and n6479_not n6480_not ; n6481
g6226 and n6478_not n6481 ; n6482
g6227 and n6215_not n6217_not ; n6483
g6228 and b[41]_not b[42]_not ; n6484
g6229 and b[41] b[42] ; n6485
g6230 and n6484_not n6485_not ; n6486
g6231 and n6483_not n6486 ; n6487
g6232 and n6483 n6486_not ; n6488
g6233 and n6487_not n6488_not ; n6489
g6234 and n269 n6489 ; n6490
g6235 and n6482 n6490_not ; n6491
g6236 and a[2] n6491_not ; n6492
g6237 and a[2] n6492_not ; n6493
g6238 and n6491_not n6492_not ; n6494
g6239 and n6493_not n6494_not ; n6495
g6240 and n6477_not n6495_not ; n6496
g6241 and n6477_not n6496_not ; n6497
g6242 and n6495_not n6496_not ; n6498
g6243 and n6497_not n6498_not ; n6499
g6244 and n6227_not n6229_not ; n6500
g6245 and n6499_not n6500_not ; n6501
g6246 and n6499 n6500 ; n6502
g6247 and n6501_not n6502_not ; f[42]
g6248 and b[43] n266 ; n6504
g6249 and b[41] n284 ; n6505
g6250 and b[42] n261 ; n6506
g6251 and n6505_not n6506_not ; n6507
g6252 and n6504_not n6507 ; n6508
g6253 and n6485_not n6487_not ; n6509
g6254 and b[42]_not b[43]_not ; n6510
g6255 and b[42] b[43] ; n6511
g6256 and n6510_not n6511_not ; n6512
g6257 and n6509_not n6512 ; n6513
g6258 and n6509 n6512_not ; n6514
g6259 and n6513_not n6514_not ; n6515
g6260 and n269 n6515 ; n6516
g6261 and n6508 n6516_not ; n6517
g6262 and a[2] n6517_not ; n6518
g6263 and a[2] n6518_not ; n6519
g6264 and n6517_not n6518_not ; n6520
g6265 and n6519_not n6520_not ; n6521
g6266 and n6470_not n6474_not ; n6522
g6267 and n6465_not n6467_not ; n6523
g6268 and b[34] n700 ; n6524
g6269 and b[32] n767 ; n6525
g6270 and b[33] n695 ; n6526
g6271 and n6525_not n6526_not ; n6527
g6272 and n6524_not n6527 ; n6528
g6273 and n703 n4466 ; n6529
g6274 and n6528 n6529_not ; n6530
g6275 and a[11] n6530_not ; n6531
g6276 and a[11] n6531_not ; n6532
g6277 and n6530_not n6531_not ; n6533
g6278 and n6532_not n6533_not ; n6534
g6279 and n6440_not n6443_not ; n6535
g6280 and n6259_not n6425_not ; n6536
g6281 and n6422_not n6536_not ; n6537
g6282 and b[28] n1302 ; n6538
g6283 and b[26] n1391 ; n6539
g6284 and b[27] n1297 ; n6540
g6285 and n6539_not n6540_not ; n6541
g6286 and n6538_not n6541 ; n6542
g6287 and n1305 n3189 ; n6543
g6288 and n6542 n6543_not ; n6544
g6289 and a[17] n6544_not ; n6545
g6290 and a[17] n6545_not ; n6546
g6291 and n6544_not n6545_not ; n6547
g6292 and n6546_not n6547_not ; n6548
g6293 and b[16] n3050 ; n6549
g6294 and b[14] n3243 ; n6550
g6295 and b[15] n3045 ; n6551
g6296 and n6550_not n6551_not ; n6552
g6297 and n6549_not n6552 ; n6553
g6298 and n1237 n3053 ; n6554
g6299 and n6553 n6554_not ; n6555
g6300 and a[29] n6555_not ; n6556
g6301 and a[29] n6556_not ; n6557
g6302 and n6555_not n6556_not ; n6558
g6303 and n6557_not n6558_not ; n6559
g6304 and n6354_not n6358_not ; n6560
g6305 and n6349_not n6351_not ; n6561
g6306 and b[7] n5035 ; n6562
g6307 and b[5] n5277 ; n6563
g6308 and b[6] n5030 ; n6564
g6309 and n6563_not n6564_not ; n6565
g6310 and n6562_not n6565 ; n6566
g6311 and n484 n5038 ; n6567
g6312 and n6566 n6567_not ; n6568
g6313 and a[38] n6568_not ; n6569
g6314 and a[38] n6569_not ; n6570
g6315 and n6568_not n6569_not ; n6571
g6316 and n6570_not n6571_not ; n6572
g6317 and n6071 n6311 ; n6573
g6318 and n6326_not n6573_not ; n6574
g6319 and b[4] n5777 ; n6575
g6320 and b[2] n6059 ; n6576
g6321 and b[3] n5772 ; n6577
g6322 and n6576_not n6577_not ; n6578
g6323 and n6575_not n6578 ; n6579
g6324 and n346 n5780 ; n6580
g6325 and n6579 n6580_not ; n6581
g6326 and a[41] n6581_not ; n6582
g6327 and a[41] n6582_not ; n6583
g6328 and n6581_not n6582_not ; n6584
g6329 and n6583_not n6584_not ; n6585
g6330 and a[44] n6311_not ; n6586
g6331 and a[42]_not a[43] ; n6587
g6332 and a[42] a[43]_not ; n6588
g6333 and n6587_not n6588_not ; n6589
g6334 and n6310 n6589_not ; n6590
g6335 and b[0] n6590 ; n6591
g6336 and a[43]_not a[44] ; n6592
g6337 and a[43] a[44]_not ; n6593
g6338 and n6592_not n6593_not ; n6594
g6339 and n6310_not n6594 ; n6595
g6340 and b[1] n6595 ; n6596
g6341 and n6591_not n6596_not ; n6597
g6342 and n6310_not n6594_not ; n6598
g6343 and n272_not n6598 ; n6599
g6344 and n6597 n6599_not ; n6600
g6345 and a[44] n6600_not ; n6601
g6346 and a[44] n6601_not ; n6602
g6347 and n6600_not n6601_not ; n6603
g6348 and n6602_not n6603_not ; n6604
g6349 and n6586 n6604_not ; n6605
g6350 and n6586_not n6604 ; n6606
g6351 and n6605_not n6606_not ; n6607
g6352 and n6585 n6607_not ; n6608
g6353 and n6585_not n6607 ; n6609
g6354 and n6608_not n6609_not ; n6610
g6355 and n6574_not n6610 ; n6611
g6356 and n6574 n6610_not ; n6612
g6357 and n6611_not n6612_not ; n6613
g6358 and n6572_not n6613 ; n6614
g6359 and n6613 n6614_not ; n6615
g6360 and n6572_not n6614_not ; n6616
g6361 and n6615_not n6616_not ; n6617
g6362 and n6329_not n6335_not ; n6618
g6363 and n6617 n6618 ; n6619
g6364 and n6617_not n6618_not ; n6620
g6365 and n6619_not n6620_not ; n6621
g6366 and b[10] n4287 ; n6622
g6367 and b[8] n4532 ; n6623
g6368 and b[9] n4282 ; n6624
g6369 and n6623_not n6624_not ; n6625
g6370 and n6622_not n6625 ; n6626
g6371 and n738 n4290 ; n6627
g6372 and n6626 n6627_not ; n6628
g6373 and a[35] n6628_not ; n6629
g6374 and a[35] n6629_not ; n6630
g6375 and n6628_not n6629_not ; n6631
g6376 and n6630_not n6631_not ; n6632
g6377 and n6621 n6632_not ; n6633
g6378 and n6621_not n6632 ; n6634
g6379 and n6561_not n6634_not ; n6635
g6380 and n6633_not n6635 ; n6636
g6381 and n6561_not n6636_not ; n6637
g6382 and n6633_not n6636_not ; n6638
g6383 and n6634_not n6638 ; n6639
g6384 and n6637_not n6639_not ; n6640
g6385 and b[13] n3638 ; n6641
g6386 and b[11] n3843 ; n6642
g6387 and b[12] n3633 ; n6643
g6388 and n6642_not n6643_not ; n6644
g6389 and n6641_not n6644 ; n6645
g6390 and n1008 n3641 ; n6646
g6391 and n6645 n6646_not ; n6647
g6392 and a[32] n6647_not ; n6648
g6393 and a[32] n6648_not ; n6649
g6394 and n6647_not n6648_not ; n6650
g6395 and n6649_not n6650_not ; n6651
g6396 and n6640 n6651 ; n6652
g6397 and n6640_not n6651_not ; n6653
g6398 and n6652_not n6653_not ; n6654
g6399 and n6560_not n6654 ; n6655
g6400 and n6560 n6654_not ; n6656
g6401 and n6655_not n6656_not ; n6657
g6402 and n6559_not n6657 ; n6658
g6403 and n6657 n6658_not ; n6659
g6404 and n6559_not n6658_not ; n6660
g6405 and n6659_not n6660_not ; n6661
g6406 and n6283_not n6376_not ; n6662
g6407 and n6373_not n6662_not ; n6663
g6408 and n6661 n6663 ; n6664
g6409 and n6661_not n6663_not ; n6665
g6410 and n6664_not n6665_not ; n6666
g6411 and b[19] n2539 ; n6667
g6412 and b[17] n2685 ; n6668
g6413 and b[18] n2534 ; n6669
g6414 and n6668_not n6669_not ; n6670
g6415 and n6667_not n6670 ; n6671
g6416 and n1708 n2542 ; n6672
g6417 and n6671 n6672_not ; n6673
g6418 and a[26] n6673_not ; n6674
g6419 and a[26] n6674_not ; n6675
g6420 and n6673_not n6674_not ; n6676
g6421 and n6675_not n6676_not ; n6677
g6422 and n6666 n6677_not ; n6678
g6423 and n6666 n6678_not ; n6679
g6424 and n6677_not n6678_not ; n6680
g6425 and n6679_not n6680_not ; n6681
g6426 and n6391_not n6394_not ; n6682
g6427 and n6681 n6682 ; n6683
g6428 and n6681_not n6682_not ; n6684
g6429 and n6683_not n6684_not ; n6685
g6430 and b[22] n2048 ; n6686
g6431 and b[20] n2198 ; n6687
g6432 and b[21] n2043 ; n6688
g6433 and n6687_not n6688_not ; n6689
g6434 and n6686_not n6689 ; n6690
g6435 and n2051 n2145 ; n6691
g6436 and n6690 n6691_not ; n6692
g6437 and a[23] n6692_not ; n6693
g6438 and a[23] n6693_not ; n6694
g6439 and n6692_not n6693_not ; n6695
g6440 and n6694_not n6695_not ; n6696
g6441 and n6685 n6696_not ; n6697
g6442 and n6685 n6697_not ; n6698
g6443 and n6696_not n6697_not ; n6699
g6444 and n6698_not n6699_not ; n6700
g6445 and n6397_not n6403_not ; n6701
g6446 and n6700 n6701 ; n6702
g6447 and n6700_not n6701_not ; n6703
g6448 and n6702_not n6703_not ; n6704
g6449 and b[25] n1627 ; n6705
g6450 and b[23] n1763 ; n6706
g6451 and b[24] n1622 ; n6707
g6452 and n6706_not n6707_not ; n6708
g6453 and n6705_not n6708 ; n6709
g6454 and n1630 n2485 ; n6710
g6455 and n6709 n6710_not ; n6711
g6456 and a[20] n6711_not ; n6712
g6457 and a[20] n6712_not ; n6713
g6458 and n6711_not n6712_not ; n6714
g6459 and n6713_not n6714_not ; n6715
g6460 and n6704 n6715_not ; n6716
g6461 and n6704 n6716_not ; n6717
g6462 and n6715_not n6716_not ; n6718
g6463 and n6717_not n6718_not ; n6719
g6464 and n6417_not n6419_not ; n6720
g6465 and n6719_not n6720_not ; n6721
g6466 and n6719 n6720 ; n6722
g6467 and n6721_not n6722_not ; n6723
g6468 and n6548_not n6723 ; n6724
g6469 and n6548_not n6724_not ; n6725
g6470 and n6723 n6724_not ; n6726
g6471 and n6725_not n6726_not ; n6727
g6472 and n6537_not n6727_not ; n6728
g6473 and n6537_not n6728_not ; n6729
g6474 and n6727_not n6728_not ; n6730
g6475 and n6729_not n6730_not ; n6731
g6476 and b[31] n951 ; n6732
g6477 and b[29] n1056 ; n6733
g6478 and b[30] n946 ; n6734
g6479 and n6733_not n6734_not ; n6735
g6480 and n6732_not n6735 ; n6736
g6481 and n954 n3796 ; n6737
g6482 and n6736 n6737_not ; n6738
g6483 and a[14] n6738_not ; n6739
g6484 and a[14] n6739_not ; n6740
g6485 and n6738_not n6739_not ; n6741
g6486 and n6740_not n6741_not ; n6742
g6487 and n6731 n6742 ; n6743
g6488 and n6731_not n6742_not ; n6744
g6489 and n6743_not n6744_not ; n6745
g6490 and n6535_not n6745 ; n6746
g6491 and n6535 n6745_not ; n6747
g6492 and n6746_not n6747_not ; n6748
g6493 and n6534_not n6748 ; n6749
g6494 and n6748 n6749_not ; n6750
g6495 and n6534_not n6749_not ; n6751
g6496 and n6750_not n6751_not ; n6752
g6497 and n6246_not n6449_not ; n6753
g6498 and n6446_not n6753_not ; n6754
g6499 and n6752 n6754 ; n6755
g6500 and n6752_not n6754_not ; n6756
g6501 and n6755_not n6756_not ; n6757
g6502 and b[37] n511 ; n6758
g6503 and b[35] n541 ; n6759
g6504 and b[36] n506 ; n6760
g6505 and n6759_not n6760_not ; n6761
g6506 and n6758_not n6761 ; n6762
g6507 and n514 n5181 ; n6763
g6508 and n6762 n6763_not ; n6764
g6509 and a[8] n6764_not ; n6765
g6510 and a[8] n6765_not ; n6766
g6511 and n6764_not n6765_not ; n6767
g6512 and n6766_not n6767_not ; n6768
g6513 and n6757 n6768_not ; n6769
g6514 and n6757_not n6768 ; n6770
g6515 and n6523_not n6770_not ; n6771
g6516 and n6769_not n6771 ; n6772
g6517 and n6523_not n6772_not ; n6773
g6518 and n6769_not n6772_not ; n6774
g6519 and n6770_not n6774 ; n6775
g6520 and n6773_not n6775_not ; n6776
g6521 and b[40] n362 ; n6777
g6522 and b[38] n403 ; n6778
g6523 and b[39] n357 ; n6779
g6524 and n6778_not n6779_not ; n6780
g6525 and n6777_not n6780 ; n6781
g6526 and n365 n5955 ; n6782
g6527 and n6781 n6782_not ; n6783
g6528 and a[5] n6783_not ; n6784
g6529 and a[5] n6784_not ; n6785
g6530 and n6783_not n6784_not ; n6786
g6531 and n6785_not n6786_not ; n6787
g6532 and n6776 n6787 ; n6788
g6533 and n6776_not n6787_not ; n6789
g6534 and n6788_not n6789_not ; n6790
g6535 and n6522_not n6790 ; n6791
g6536 and n6522 n6790_not ; n6792
g6537 and n6791_not n6792_not ; n6793
g6538 and n6521_not n6793 ; n6794
g6539 and n6793 n6794_not ; n6795
g6540 and n6521_not n6794_not ; n6796
g6541 and n6795_not n6796_not ; n6797
g6542 and n6496_not n6501_not ; n6798
g6543 and n6797_not n6798_not ; n6799
g6544 and n6797 n6798 ; n6800
g6545 and n6799_not n6800_not ; f[43]
g6546 and n6794_not n6799_not ; n6802
g6547 and n6789_not n6791_not ; n6803
g6548 and b[41] n362 ; n6804
g6549 and b[39] n403 ; n6805
g6550 and b[40] n357 ; n6806
g6551 and n6805_not n6806_not ; n6807
g6552 and n6804_not n6807 ; n6808
g6553 and n365 n6219 ; n6809
g6554 and n6808 n6809_not ; n6810
g6555 and a[5] n6810_not ; n6811
g6556 and a[5] n6811_not ; n6812
g6557 and n6810_not n6811_not ; n6813
g6558 and n6812_not n6813_not ; n6814
g6559 and b[35] n700 ; n6815
g6560 and b[33] n767 ; n6816
g6561 and b[34] n695 ; n6817
g6562 and n6816_not n6817_not ; n6818
g6563 and n6815_not n6818 ; n6819
g6564 and n703 n4696 ; n6820
g6565 and n6819 n6820_not ; n6821
g6566 and a[11] n6821_not ; n6822
g6567 and a[11] n6822_not ; n6823
g6568 and n6821_not n6822_not ; n6824
g6569 and n6823_not n6824_not ; n6825
g6570 and n6744_not n6746_not ; n6826
g6571 and b[32] n951 ; n6827
g6572 and b[30] n1056 ; n6828
g6573 and b[31] n946 ; n6829
g6574 and n6828_not n6829_not ; n6830
g6575 and n6827_not n6830 ; n6831
g6576 and n954 n4013 ; n6832
g6577 and n6831 n6832_not ; n6833
g6578 and a[14] n6833_not ; n6834
g6579 and a[14] n6834_not ; n6835
g6580 and n6833_not n6834_not ; n6836
g6581 and n6835_not n6836_not ; n6837
g6582 and n6724_not n6728_not ; n6838
g6583 and b[29] n1302 ; n6839
g6584 and b[27] n1391 ; n6840
g6585 and b[28] n1297 ; n6841
g6586 and n6840_not n6841_not ; n6842
g6587 and n6839_not n6842 ; n6843
g6588 and n1305 n3383 ; n6844
g6589 and n6843 n6844_not ; n6845
g6590 and a[17] n6845_not ; n6846
g6591 and a[17] n6846_not ; n6847
g6592 and n6845_not n6846_not ; n6848
g6593 and n6847_not n6848_not ; n6849
g6594 and n6716_not n6721_not ; n6850
g6595 and n6697_not n6703_not ; n6851
g6596 and b[20] n2539 ; n6852
g6597 and b[18] n2685 ; n6853
g6598 and b[19] n2534 ; n6854
g6599 and n6853_not n6854_not ; n6855
g6600 and n6852_not n6855 ; n6856
g6601 and n1846 n2542 ; n6857
g6602 and n6856 n6857_not ; n6858
g6603 and a[26] n6858_not ; n6859
g6604 and a[26] n6859_not ; n6860
g6605 and n6858_not n6859_not ; n6861
g6606 and n6860_not n6861_not ; n6862
g6607 and n6658_not n6665_not ; n6863
g6608 and b[17] n3050 ; n6864
g6609 and b[15] n3243 ; n6865
g6610 and b[16] n3045 ; n6866
g6611 and n6865_not n6866_not ; n6867
g6612 and n6864_not n6867 ; n6868
g6613 and n1356 n3053 ; n6869
g6614 and n6868 n6869_not ; n6870
g6615 and a[29] n6870_not ; n6871
g6616 and a[29] n6871_not ; n6872
g6617 and n6870_not n6871_not ; n6873
g6618 and n6872_not n6873_not ; n6874
g6619 and n6653_not n6655_not ; n6875
g6620 and b[14] n3638 ; n6876
g6621 and b[12] n3843 ; n6877
g6622 and b[13] n3633 ; n6878
g6623 and n6877_not n6878_not ; n6879
g6624 and n6876_not n6879 ; n6880
g6625 and n1034 n3641 ; n6881
g6626 and n6880 n6881_not ; n6882
g6627 and a[32] n6882_not ; n6883
g6628 and a[32] n6883_not ; n6884
g6629 and n6882_not n6883_not ; n6885
g6630 and n6884_not n6885_not ; n6886
g6631 and n6614_not n6620_not ; n6887
g6632 and b[8] n5035 ; n6888
g6633 and b[6] n5277 ; n6889
g6634 and b[7] n5030 ; n6890
g6635 and n6889_not n6890_not ; n6891
g6636 and n6888_not n6891 ; n6892
g6637 and n585 n5038 ; n6893
g6638 and n6892 n6893_not ; n6894
g6639 and a[38] n6894_not ; n6895
g6640 and a[38] n6895_not ; n6896
g6641 and n6894_not n6895_not ; n6897
g6642 and n6896_not n6897_not ; n6898
g6643 and n6609_not n6611_not ; n6899
g6644 and b[2] n6595 ; n6900
g6645 and n6310 n6594_not ; n6901
g6646 and n6589 n6901 ; n6902
g6647 and b[0] n6902 ; n6903
g6648 and b[1] n6590 ; n6904
g6649 and n6903_not n6904_not ; n6905
g6650 and n6900_not n6905 ; n6906
g6651 and n296 n6598 ; n6907
g6652 and n6906 n6907_not ; n6908
g6653 and a[44] n6908_not ; n6909
g6654 and a[44] n6909_not ; n6910
g6655 and n6908_not n6909_not ; n6911
g6656 and n6910_not n6911_not ; n6912
g6657 and n6605_not n6912 ; n6913
g6658 and n6605 n6912_not ; n6914
g6659 and n6913_not n6914_not ; n6915
g6660 and b[5] n5777 ; n6916
g6661 and b[3] n6059 ; n6917
g6662 and b[4] n5772 ; n6918
g6663 and n6917_not n6918_not ; n6919
g6664 and n6916_not n6919 ; n6920
g6665 and n394 n5780 ; n6921
g6666 and n6920 n6921_not ; n6922
g6667 and a[41] n6922_not ; n6923
g6668 and a[41] n6923_not ; n6924
g6669 and n6922_not n6923_not ; n6925
g6670 and n6924_not n6925_not ; n6926
g6671 and n6915 n6926_not ; n6927
g6672 and n6915 n6927_not ; n6928
g6673 and n6926_not n6927_not ; n6929
g6674 and n6928_not n6929_not ; n6930
g6675 and n6899_not n6930_not ; n6931
g6676 and n6899 n6930 ; n6932
g6677 and n6931_not n6932_not ; n6933
g6678 and n6898_not n6933 ; n6934
g6679 and n6898_not n6934_not ; n6935
g6680 and n6933 n6934_not ; n6936
g6681 and n6935_not n6936_not ; n6937
g6682 and n6887_not n6937_not ; n6938
g6683 and n6887_not n6938_not ; n6939
g6684 and n6937_not n6938_not ; n6940
g6685 and n6939_not n6940_not ; n6941
g6686 and b[11] n4287 ; n6942
g6687 and b[9] n4532 ; n6943
g6688 and b[10] n4282 ; n6944
g6689 and n6943_not n6944_not ; n6945
g6690 and n6942_not n6945 ; n6946
g6691 and n818 n4290 ; n6947
g6692 and n6946 n6947_not ; n6948
g6693 and a[35] n6948_not ; n6949
g6694 and a[35] n6949_not ; n6950
g6695 and n6948_not n6949_not ; n6951
g6696 and n6950_not n6951_not ; n6952
g6697 and n6941 n6952 ; n6953
g6698 and n6941_not n6952_not ; n6954
g6699 and n6953_not n6954_not ; n6955
g6700 and n6638_not n6955 ; n6956
g6701 and n6638 n6955_not ; n6957
g6702 and n6956_not n6957_not ; n6958
g6703 and n6886 n6958_not ; n6959
g6704 and n6886_not n6958 ; n6960
g6705 and n6959_not n6960_not ; n6961
g6706 and n6875_not n6961 ; n6962
g6707 and n6875 n6961_not ; n6963
g6708 and n6962_not n6963_not ; n6964
g6709 and n6874 n6964_not ; n6965
g6710 and n6874_not n6964 ; n6966
g6711 and n6965_not n6966_not ; n6967
g6712 and n6863_not n6967 ; n6968
g6713 and n6863 n6967_not ; n6969
g6714 and n6968_not n6969_not ; n6970
g6715 and n6862_not n6970 ; n6971
g6716 and n6970 n6971_not ; n6972
g6717 and n6862_not n6971_not ; n6973
g6718 and n6972_not n6973_not ; n6974
g6719 and n6678_not n6684_not ; n6975
g6720 and n6974 n6975 ; n6976
g6721 and n6974_not n6975_not ; n6977
g6722 and n6976_not n6977_not ; n6978
g6723 and b[23] n2048 ; n6979
g6724 and b[21] n2198 ; n6980
g6725 and b[22] n2043 ; n6981
g6726 and n6980_not n6981_not ; n6982
g6727 and n6979_not n6982 ; n6983
g6728 and n2051 n2300 ; n6984
g6729 and n6983 n6984_not ; n6985
g6730 and a[23] n6985_not ; n6986
g6731 and a[23] n6986_not ; n6987
g6732 and n6985_not n6986_not ; n6988
g6733 and n6987_not n6988_not ; n6989
g6734 and n6978 n6989_not ; n6990
g6735 and n6978_not n6989 ; n6991
g6736 and n6851_not n6991_not ; n6992
g6737 and n6990_not n6992 ; n6993
g6738 and n6851_not n6993_not ; n6994
g6739 and n6990_not n6993_not ; n6995
g6740 and n6991_not n6995 ; n6996
g6741 and n6994_not n6996_not ; n6997
g6742 and b[26] n1627 ; n6998
g6743 and b[24] n1763 ; n6999
g6744 and b[25] n1622 ; n7000
g6745 and n6999_not n7000_not ; n7001
g6746 and n6998_not n7001 ; n7002
g6747 and n1630 n2813 ; n7003
g6748 and n7002 n7003_not ; n7004
g6749 and a[20] n7004_not ; n7005
g6750 and a[20] n7005_not ; n7006
g6751 and n7004_not n7005_not ; n7007
g6752 and n7006_not n7007_not ; n7008
g6753 and n6997 n7008 ; n7009
g6754 and n6997_not n7008_not ; n7010
g6755 and n7009_not n7010_not ; n7011
g6756 and n6850_not n7011 ; n7012
g6757 and n6850 n7011_not ; n7013
g6758 and n7012_not n7013_not ; n7014
g6759 and n6849 n7014_not ; n7015
g6760 and n6849_not n7014 ; n7016
g6761 and n7015_not n7016_not ; n7017
g6762 and n6838_not n7017 ; n7018
g6763 and n6838 n7017_not ; n7019
g6764 and n7018_not n7019_not ; n7020
g6765 and n6837 n7020_not ; n7021
g6766 and n6837_not n7020 ; n7022
g6767 and n7021_not n7022_not ; n7023
g6768 and n6826_not n7023 ; n7024
g6769 and n6826 n7023_not ; n7025
g6770 and n7024_not n7025_not ; n7026
g6771 and n6825_not n7026 ; n7027
g6772 and n7026 n7027_not ; n7028
g6773 and n6825_not n7027_not ; n7029
g6774 and n7028_not n7029_not ; n7030
g6775 and n6749_not n6756_not ; n7031
g6776 and n7030 n7031 ; n7032
g6777 and n7030_not n7031_not ; n7033
g6778 and n7032_not n7033_not ; n7034
g6779 and b[38] n511 ; n7035
g6780 and b[36] n541 ; n7036
g6781 and b[37] n506 ; n7037
g6782 and n7036_not n7037_not ; n7038
g6783 and n7035_not n7038 ; n7039
g6784 and n514 n5205 ; n7040
g6785 and n7039 n7040_not ; n7041
g6786 and a[8] n7041_not ; n7042
g6787 and a[8] n7042_not ; n7043
g6788 and n7041_not n7042_not ; n7044
g6789 and n7043_not n7044_not ; n7045
g6790 and n7034 n7045_not ; n7046
g6791 and n7034 n7046_not ; n7047
g6792 and n7045_not n7046_not ; n7048
g6793 and n7047_not n7048_not ; n7049
g6794 and n6774_not n7049_not ; n7050
g6795 and n6774 n7049 ; n7051
g6796 and n7050_not n7051_not ; n7052
g6797 and n6814_not n7052 ; n7053
g6798 and n6814_not n7053_not ; n7054
g6799 and n7052 n7053_not ; n7055
g6800 and n7054_not n7055_not ; n7056
g6801 and n6803_not n7056_not ; n7057
g6802 and n6803_not n7057_not ; n7058
g6803 and n7056_not n7057_not ; n7059
g6804 and n7058_not n7059_not ; n7060
g6805 and b[44] n266 ; n7061
g6806 and b[42] n284 ; n7062
g6807 and b[43] n261 ; n7063
g6808 and n7062_not n7063_not ; n7064
g6809 and n7061_not n7064 ; n7065
g6810 and n6511_not n6513_not ; n7066
g6811 and b[43]_not b[44]_not ; n7067
g6812 and b[43] b[44] ; n7068
g6813 and n7067_not n7068_not ; n7069
g6814 and n7066_not n7069 ; n7070
g6815 and n7066 n7069_not ; n7071
g6816 and n7070_not n7071_not ; n7072
g6817 and n269 n7072 ; n7073
g6818 and n7065 n7073_not ; n7074
g6819 and a[2] n7074_not ; n7075
g6820 and a[2] n7075_not ; n7076
g6821 and n7074_not n7075_not ; n7077
g6822 and n7076_not n7077_not ; n7078
g6823 and n7060_not n7078 ; n7079
g6824 and n7060 n7078_not ; n7080
g6825 and n7079_not n7080_not ; n7081
g6826 and n6802_not n7081_not ; n7082
g6827 and n6802 n7081 ; n7083
g6828 and n7082_not n7083_not ; f[44]
g6829 and n7060_not n7078_not ; n7085
g6830 and n7082_not n7085_not ; n7086
g6831 and n7027_not n7033_not ; n7087
g6832 and n7022_not n7024_not ; n7088
g6833 and b[33] n951 ; n7089
g6834 and b[31] n1056 ; n7090
g6835 and b[32] n946 ; n7091
g6836 and n7090_not n7091_not ; n7092
g6837 and n7089_not n7092 ; n7093
g6838 and n954 n4223 ; n7094
g6839 and n7093 n7094_not ; n7095
g6840 and a[14] n7095_not ; n7096
g6841 and a[14] n7096_not ; n7097
g6842 and n7095_not n7096_not ; n7098
g6843 and n7097_not n7098_not ; n7099
g6844 and n7016_not n7018_not ; n7100
g6845 and n7010_not n7012_not ; n7101
g6846 and b[27] n1627 ; n7102
g6847 and b[25] n1763 ; n7103
g6848 and b[26] n1622 ; n7104
g6849 and n7103_not n7104_not ; n7105
g6850 and n7102_not n7105 ; n7106
g6851 and n1630 n2990 ; n7107
g6852 and n7106 n7107_not ; n7108
g6853 and a[20] n7108_not ; n7109
g6854 and a[20] n7109_not ; n7110
g6855 and n7108_not n7109_not ; n7111
g6856 and n7110_not n7111_not ; n7112
g6857 and b[21] n2539 ; n7113
g6858 and b[19] n2685 ; n7114
g6859 and b[20] n2534 ; n7115
g6860 and n7114_not n7115_not ; n7116
g6861 and n7113_not n7116 ; n7117
g6862 and n1984 n2542 ; n7118
g6863 and n7117 n7118_not ; n7119
g6864 and a[26] n7119_not ; n7120
g6865 and a[26] n7120_not ; n7121
g6866 and n7119_not n7120_not ; n7122
g6867 and n7121_not n7122_not ; n7123
g6868 and n6966_not n6968_not ; n7124
g6869 and n6960_not n6962_not ; n7125
g6870 and n6954_not n6956_not ; n7126
g6871 and b[12] n4287 ; n7127
g6872 and b[10] n4532 ; n7128
g6873 and b[11] n4282 ; n7129
g6874 and n7128_not n7129_not ; n7130
g6875 and n7127_not n7130 ; n7131
g6876 and n842 n4290 ; n7132
g6877 and n7131 n7132_not ; n7133
g6878 and a[35] n7133_not ; n7134
g6879 and a[35] n7134_not ; n7135
g6880 and n7133_not n7134_not ; n7136
g6881 and n7135_not n7136_not ; n7137
g6882 and n6934_not n6938_not ; n7138
g6883 and b[6] n5777 ; n7139
g6884 and b[4] n6059 ; n7140
g6885 and b[5] n5772 ; n7141
g6886 and n7140_not n7141_not ; n7142
g6887 and n7139_not n7142 ; n7143
g6888 and n459 n5780 ; n7144
g6889 and n7143 n7144_not ; n7145
g6890 and a[41] n7145_not ; n7146
g6891 and a[41] n7146_not ; n7147
g6892 and n7145_not n7146_not ; n7148
g6893 and n7147_not n7148_not ; n7149
g6894 and a[44] a[45]_not ; n7150
g6895 and a[44]_not a[45] ; n7151
g6896 and n7150_not n7151_not ; n7152
g6897 and b[0] n7152_not ; n7153
g6898 and n6914_not n7153 ; n7154
g6899 and n6914 n7153_not ; n7155
g6900 and n7154_not n7155_not ; n7156
g6901 and b[3] n6595 ; n7157
g6902 and b[1] n6902 ; n7158
g6903 and b[2] n6590 ; n7159
g6904 and n7158_not n7159_not ; n7160
g6905 and n7157_not n7160 ; n7161
g6906 and n318 n6598 ; n7162
g6907 and n7161 n7162_not ; n7163
g6908 and a[44] n7163_not ; n7164
g6909 and a[44] n7164_not ; n7165
g6910 and n7163_not n7164_not ; n7166
g6911 and n7165_not n7166_not ; n7167
g6912 and n7156_not n7167_not ; n7168
g6913 and n7156 n7167 ; n7169
g6914 and n7168_not n7169_not ; n7170
g6915 and n7149_not n7170 ; n7171
g6916 and n7170 n7171_not ; n7172
g6917 and n7149_not n7171_not ; n7173
g6918 and n7172_not n7173_not ; n7174
g6919 and n6927_not n6931_not ; n7175
g6920 and n7174 n7175 ; n7176
g6921 and n7174_not n7175_not ; n7177
g6922 and n7176_not n7177_not ; n7178
g6923 and b[9] n5035 ; n7179
g6924 and b[7] n5277 ; n7180
g6925 and b[8] n5030 ; n7181
g6926 and n7180_not n7181_not ; n7182
g6927 and n7179_not n7182 ; n7183
g6928 and n651 n5038 ; n7184
g6929 and n7183 n7184_not ; n7185
g6930 and a[38] n7185_not ; n7186
g6931 and a[38] n7186_not ; n7187
g6932 and n7185_not n7186_not ; n7188
g6933 and n7187_not n7188_not ; n7189
g6934 and n7178_not n7189 ; n7190
g6935 and n7178 n7189_not ; n7191
g6936 and n7190_not n7191_not ; n7192
g6937 and n7138_not n7192 ; n7193
g6938 and n7138 n7192_not ; n7194
g6939 and n7193_not n7194_not ; n7195
g6940 and n7137_not n7195 ; n7196
g6941 and n7137_not n7196_not ; n7197
g6942 and n7195 n7196_not ; n7198
g6943 and n7197_not n7198_not ; n7199
g6944 and n7126_not n7199_not ; n7200
g6945 and n7126_not n7200_not ; n7201
g6946 and n7199_not n7200_not ; n7202
g6947 and n7201_not n7202_not ; n7203
g6948 and b[15] n3638 ; n7204
g6949 and b[13] n3843 ; n7205
g6950 and b[14] n3633 ; n7206
g6951 and n7205_not n7206_not ; n7207
g6952 and n7204_not n7207 ; n7208
g6953 and n1131 n3641 ; n7209
g6954 and n7208 n7209_not ; n7210
g6955 and a[32] n7210_not ; n7211
g6956 and a[32] n7211_not ; n7212
g6957 and n7210_not n7211_not ; n7213
g6958 and n7212_not n7213_not ; n7214
g6959 and n7203_not n7214_not ; n7215
g6960 and n7203_not n7215_not ; n7216
g6961 and n7214_not n7215_not ; n7217
g6962 and n7216_not n7217_not ; n7218
g6963 and n7125_not n7218 ; n7219
g6964 and n7125 n7218_not ; n7220
g6965 and n7219_not n7220_not ; n7221
g6966 and b[18] n3050 ; n7222
g6967 and b[16] n3243 ; n7223
g6968 and b[17] n3045 ; n7224
g6969 and n7223_not n7224_not ; n7225
g6970 and n7222_not n7225 ; n7226
g6971 and n1566 n3053 ; n7227
g6972 and n7226 n7227_not ; n7228
g6973 and a[29] n7228_not ; n7229
g6974 and a[29] n7229_not ; n7230
g6975 and n7228_not n7229_not ; n7231
g6976 and n7230_not n7231_not ; n7232
g6977 and n7221_not n7232_not ; n7233
g6978 and n7221 n7232 ; n7234
g6979 and n7233_not n7234_not ; n7235
g6980 and n7124_not n7235 ; n7236
g6981 and n7124 n7235_not ; n7237
g6982 and n7236_not n7237_not ; n7238
g6983 and n7123_not n7238 ; n7239
g6984 and n7238 n7239_not ; n7240
g6985 and n7123_not n7239_not ; n7241
g6986 and n7240_not n7241_not ; n7242
g6987 and n6971_not n6977_not ; n7243
g6988 and n7242 n7243 ; n7244
g6989 and n7242_not n7243_not ; n7245
g6990 and n7244_not n7245_not ; n7246
g6991 and b[24] n2048 ; n7247
g6992 and b[22] n2198 ; n7248
g6993 and b[23] n2043 ; n7249
g6994 and n7248_not n7249_not ; n7250
g6995 and n7247_not n7250 ; n7251
g6996 and n2051 n2458 ; n7252
g6997 and n7251 n7252_not ; n7253
g6998 and a[23] n7253_not ; n7254
g6999 and a[23] n7254_not ; n7255
g7000 and n7253_not n7254_not ; n7256
g7001 and n7255_not n7256_not ; n7257
g7002 and n7246_not n7257 ; n7258
g7003 and n7246 n7257_not ; n7259
g7004 and n7258_not n7259_not ; n7260
g7005 and n6995_not n7260 ; n7261
g7006 and n6995 n7260_not ; n7262
g7007 and n7261_not n7262_not ; n7263
g7008 and n7112_not n7263 ; n7264
g7009 and n7263 n7264_not ; n7265
g7010 and n7112_not n7264_not ; n7266
g7011 and n7265_not n7266_not ; n7267
g7012 and n7101_not n7267 ; n7268
g7013 and n7101 n7267_not ; n7269
g7014 and n7268_not n7269_not ; n7270
g7015 and b[30] n1302 ; n7271
g7016 and b[28] n1391 ; n7272
g7017 and b[29] n1297 ; n7273
g7018 and n7272_not n7273_not ; n7274
g7019 and n7271_not n7274 ; n7275
g7020 and n1305 n3577 ; n7276
g7021 and n7275 n7276_not ; n7277
g7022 and a[17] n7277_not ; n7278
g7023 and a[17] n7278_not ; n7279
g7024 and n7277_not n7278_not ; n7280
g7025 and n7279_not n7280_not ; n7281
g7026 and n7270_not n7281_not ; n7282
g7027 and n7270 n7281 ; n7283
g7028 and n7282_not n7283_not ; n7284
g7029 and n7100_not n7284 ; n7285
g7030 and n7100 n7284_not ; n7286
g7031 and n7285_not n7286_not ; n7287
g7032 and n7099_not n7287 ; n7288
g7033 and n7287 n7288_not ; n7289
g7034 and n7099_not n7288_not ; n7290
g7035 and n7289_not n7290_not ; n7291
g7036 and n7088_not n7291 ; n7292
g7037 and n7088 n7291_not ; n7293
g7038 and n7292_not n7293_not ; n7294
g7039 and b[36] n700 ; n7295
g7040 and b[34] n767 ; n7296
g7041 and b[35] n695 ; n7297
g7042 and n7296_not n7297_not ; n7298
g7043 and n7295_not n7298 ; n7299
g7044 and n703 n4922 ; n7300
g7045 and n7299 n7300_not ; n7301
g7046 and a[11] n7301_not ; n7302
g7047 and a[11] n7302_not ; n7303
g7048 and n7301_not n7302_not ; n7304
g7049 and n7303_not n7304_not ; n7305
g7050 and n7294_not n7305_not ; n7306
g7051 and n7294 n7305 ; n7307
g7052 and n7306_not n7307_not ; n7308
g7053 and n7087 n7308_not ; n7309
g7054 and n7087_not n7308 ; n7310
g7055 and n7309_not n7310_not ; n7311
g7056 and b[39] n511 ; n7312
g7057 and b[37] n541 ; n7313
g7058 and b[38] n506 ; n7314
g7059 and n7313_not n7314_not ; n7315
g7060 and n7312_not n7315 ; n7316
g7061 and n514 n5451 ; n7317
g7062 and n7316 n7317_not ; n7318
g7063 and a[8] n7318_not ; n7319
g7064 and a[8] n7319_not ; n7320
g7065 and n7318_not n7319_not ; n7321
g7066 and n7320_not n7321_not ; n7322
g7067 and n7311 n7322_not ; n7323
g7068 and n7311 n7323_not ; n7324
g7069 and n7322_not n7323_not ; n7325
g7070 and n7324_not n7325_not ; n7326
g7071 and n7046_not n7050_not ; n7327
g7072 and n7326 n7327 ; n7328
g7073 and n7326_not n7327_not ; n7329
g7074 and n7328_not n7329_not ; n7330
g7075 and b[42] n362 ; n7331
g7076 and b[40] n403 ; n7332
g7077 and b[41] n357 ; n7333
g7078 and n7332_not n7333_not ; n7334
g7079 and n7331_not n7334 ; n7335
g7080 and n365 n6489 ; n7336
g7081 and n7335 n7336_not ; n7337
g7082 and a[5] n7337_not ; n7338
g7083 and a[5] n7338_not ; n7339
g7084 and n7337_not n7338_not ; n7340
g7085 and n7339_not n7340_not ; n7341
g7086 and n7330 n7341_not ; n7342
g7087 and n7330 n7342_not ; n7343
g7088 and n7341_not n7342_not ; n7344
g7089 and n7343_not n7344_not ; n7345
g7090 and n7053_not n7057_not ; n7346
g7091 and n7345 n7346 ; n7347
g7092 and n7345_not n7346_not ; n7348
g7093 and n7347_not n7348_not ; n7349
g7094 and b[45] n266 ; n7350
g7095 and b[43] n284 ; n7351
g7096 and b[44] n261 ; n7352
g7097 and n7351_not n7352_not ; n7353
g7098 and n7350_not n7353 ; n7354
g7099 and n7068_not n7070_not ; n7355
g7100 and b[44]_not b[45]_not ; n7356
g7101 and b[44] b[45] ; n7357
g7102 and n7356_not n7357_not ; n7358
g7103 and n7355_not n7358 ; n7359
g7104 and n7355 n7358_not ; n7360
g7105 and n7359_not n7360_not ; n7361
g7106 and n269 n7361 ; n7362
g7107 and n7354 n7362_not ; n7363
g7108 and a[2] n7363_not ; n7364
g7109 and a[2] n7364_not ; n7365
g7110 and n7363_not n7364_not ; n7366
g7111 and n7365_not n7366_not ; n7367
g7112 and n7349_not n7367 ; n7368
g7113 and n7349 n7367_not ; n7369
g7114 and n7368_not n7369_not ; n7370
g7115 and n7086_not n7370 ; n7371
g7116 and n7086 n7370_not ; n7372
g7117 and n7371_not n7372_not ; f[45]
g7118 and n7323_not n7329_not ; n7374
g7119 and b[34] n951 ; n7375
g7120 and b[32] n1056 ; n7376
g7121 and b[33] n946 ; n7377
g7122 and n7376_not n7377_not ; n7378
g7123 and n7375_not n7378 ; n7379
g7124 and n954 n4466 ; n7380
g7125 and n7379 n7380_not ; n7381
g7126 and a[14] n7381_not ; n7382
g7127 and a[14] n7382_not ; n7383
g7128 and n7381_not n7382_not ; n7384
g7129 and n7383_not n7384_not ; n7385
g7130 and n7282_not n7285_not ; n7386
g7131 and n7101_not n7267_not ; n7387
g7132 and n7264_not n7387_not ; n7388
g7133 and b[28] n1627 ; n7389
g7134 and b[26] n1763 ; n7390
g7135 and b[27] n1622 ; n7391
g7136 and n7390_not n7391_not ; n7392
g7137 and n7389_not n7392 ; n7393
g7138 and n1630 n3189 ; n7394
g7139 and n7393 n7394_not ; n7395
g7140 and a[20] n7395_not ; n7396
g7141 and a[20] n7396_not ; n7397
g7142 and n7395_not n7396_not ; n7398
g7143 and n7397_not n7398_not ; n7399
g7144 and b[16] n3638 ; n7400
g7145 and b[14] n3843 ; n7401
g7146 and b[15] n3633 ; n7402
g7147 and n7401_not n7402_not ; n7403
g7148 and n7400_not n7403 ; n7404
g7149 and n1237 n3641 ; n7405
g7150 and n7404 n7405_not ; n7406
g7151 and a[32] n7406_not ; n7407
g7152 and a[32] n7407_not ; n7408
g7153 and n7406_not n7407_not ; n7409
g7154 and n7408_not n7409_not ; n7410
g7155 and n7196_not n7200_not ; n7411
g7156 and n7191_not n7193_not ; n7412
g7157 and b[7] n5777 ; n7413
g7158 and b[5] n6059 ; n7414
g7159 and b[6] n5772 ; n7415
g7160 and n7414_not n7415_not ; n7416
g7161 and n7413_not n7416 ; n7417
g7162 and n484 n5780 ; n7418
g7163 and n7417 n7418_not ; n7419
g7164 and a[41] n7419_not ; n7420
g7165 and a[41] n7420_not ; n7421
g7166 and n7419_not n7420_not ; n7422
g7167 and n7421_not n7422_not ; n7423
g7168 and n6914 n7153 ; n7424
g7169 and n7168_not n7424_not ; n7425
g7170 and b[4] n6595 ; n7426
g7171 and b[2] n6902 ; n7427
g7172 and b[3] n6590 ; n7428
g7173 and n7427_not n7428_not ; n7429
g7174 and n7426_not n7429 ; n7430
g7175 and n346 n6598 ; n7431
g7176 and n7430 n7431_not ; n7432
g7177 and a[44] n7432_not ; n7433
g7178 and a[44] n7433_not ; n7434
g7179 and n7432_not n7433_not ; n7435
g7180 and n7434_not n7435_not ; n7436
g7181 and a[47] n7153_not ; n7437
g7182 and a[45]_not a[46] ; n7438
g7183 and a[45] a[46]_not ; n7439
g7184 and n7438_not n7439_not ; n7440
g7185 and n7152 n7440_not ; n7441
g7186 and b[0] n7441 ; n7442
g7187 and a[46]_not a[47] ; n7443
g7188 and a[46] a[47]_not ; n7444
g7189 and n7443_not n7444_not ; n7445
g7190 and n7152_not n7445 ; n7446
g7191 and b[1] n7446 ; n7447
g7192 and n7442_not n7447_not ; n7448
g7193 and n7152_not n7445_not ; n7449
g7194 and n272_not n7449 ; n7450
g7195 and n7448 n7450_not ; n7451
g7196 and a[47] n7451_not ; n7452
g7197 and a[47] n7452_not ; n7453
g7198 and n7451_not n7452_not ; n7454
g7199 and n7453_not n7454_not ; n7455
g7200 and n7437 n7455_not ; n7456
g7201 and n7437_not n7455 ; n7457
g7202 and n7456_not n7457_not ; n7458
g7203 and n7436 n7458_not ; n7459
g7204 and n7436_not n7458 ; n7460
g7205 and n7459_not n7460_not ; n7461
g7206 and n7425_not n7461 ; n7462
g7207 and n7425 n7461_not ; n7463
g7208 and n7462_not n7463_not ; n7464
g7209 and n7423_not n7464 ; n7465
g7210 and n7464 n7465_not ; n7466
g7211 and n7423_not n7465_not ; n7467
g7212 and n7466_not n7467_not ; n7468
g7213 and n7171_not n7177_not ; n7469
g7214 and n7468 n7469 ; n7470
g7215 and n7468_not n7469_not ; n7471
g7216 and n7470_not n7471_not ; n7472
g7217 and b[10] n5035 ; n7473
g7218 and b[8] n5277 ; n7474
g7219 and b[9] n5030 ; n7475
g7220 and n7474_not n7475_not ; n7476
g7221 and n7473_not n7476 ; n7477
g7222 and n738 n5038 ; n7478
g7223 and n7477 n7478_not ; n7479
g7224 and a[38] n7479_not ; n7480
g7225 and a[38] n7480_not ; n7481
g7226 and n7479_not n7480_not ; n7482
g7227 and n7481_not n7482_not ; n7483
g7228 and n7472 n7483_not ; n7484
g7229 and n7472_not n7483 ; n7485
g7230 and n7412_not n7485_not ; n7486
g7231 and n7484_not n7486 ; n7487
g7232 and n7412_not n7487_not ; n7488
g7233 and n7484_not n7487_not ; n7489
g7234 and n7485_not n7489 ; n7490
g7235 and n7488_not n7490_not ; n7491
g7236 and b[13] n4287 ; n7492
g7237 and b[11] n4532 ; n7493
g7238 and b[12] n4282 ; n7494
g7239 and n7493_not n7494_not ; n7495
g7240 and n7492_not n7495 ; n7496
g7241 and n1008 n4290 ; n7497
g7242 and n7496 n7497_not ; n7498
g7243 and a[35] n7498_not ; n7499
g7244 and a[35] n7499_not ; n7500
g7245 and n7498_not n7499_not ; n7501
g7246 and n7500_not n7501_not ; n7502
g7247 and n7491 n7502 ; n7503
g7248 and n7491_not n7502_not ; n7504
g7249 and n7503_not n7504_not ; n7505
g7250 and n7411_not n7505 ; n7506
g7251 and n7411 n7505_not ; n7507
g7252 and n7506_not n7507_not ; n7508
g7253 and n7410_not n7508 ; n7509
g7254 and n7508 n7509_not ; n7510
g7255 and n7410_not n7509_not ; n7511
g7256 and n7510_not n7511_not ; n7512
g7257 and n7125_not n7218_not ; n7513
g7258 and n7215_not n7513_not ; n7514
g7259 and n7512 n7514 ; n7515
g7260 and n7512_not n7514_not ; n7516
g7261 and n7515_not n7516_not ; n7517
g7262 and b[19] n3050 ; n7518
g7263 and b[17] n3243 ; n7519
g7264 and b[18] n3045 ; n7520
g7265 and n7519_not n7520_not ; n7521
g7266 and n7518_not n7521 ; n7522
g7267 and n1708 n3053 ; n7523
g7268 and n7522 n7523_not ; n7524
g7269 and a[29] n7524_not ; n7525
g7270 and a[29] n7525_not ; n7526
g7271 and n7524_not n7525_not ; n7527
g7272 and n7526_not n7527_not ; n7528
g7273 and n7517 n7528_not ; n7529
g7274 and n7517 n7529_not ; n7530
g7275 and n7528_not n7529_not ; n7531
g7276 and n7530_not n7531_not ; n7532
g7277 and n7233_not n7236_not ; n7533
g7278 and n7532 n7533 ; n7534
g7279 and n7532_not n7533_not ; n7535
g7280 and n7534_not n7535_not ; n7536
g7281 and b[22] n2539 ; n7537
g7282 and b[20] n2685 ; n7538
g7283 and b[21] n2534 ; n7539
g7284 and n7538_not n7539_not ; n7540
g7285 and n7537_not n7540 ; n7541
g7286 and n2145 n2542 ; n7542
g7287 and n7541 n7542_not ; n7543
g7288 and a[26] n7543_not ; n7544
g7289 and a[26] n7544_not ; n7545
g7290 and n7543_not n7544_not ; n7546
g7291 and n7545_not n7546_not ; n7547
g7292 and n7536 n7547_not ; n7548
g7293 and n7536 n7548_not ; n7549
g7294 and n7547_not n7548_not ; n7550
g7295 and n7549_not n7550_not ; n7551
g7296 and n7239_not n7245_not ; n7552
g7297 and n7551 n7552 ; n7553
g7298 and n7551_not n7552_not ; n7554
g7299 and n7553_not n7554_not ; n7555
g7300 and b[25] n2048 ; n7556
g7301 and b[23] n2198 ; n7557
g7302 and b[24] n2043 ; n7558
g7303 and n7557_not n7558_not ; n7559
g7304 and n7556_not n7559 ; n7560
g7305 and n2051 n2485 ; n7561
g7306 and n7560 n7561_not ; n7562
g7307 and a[23] n7562_not ; n7563
g7308 and a[23] n7563_not ; n7564
g7309 and n7562_not n7563_not ; n7565
g7310 and n7564_not n7565_not ; n7566
g7311 and n7555 n7566_not ; n7567
g7312 and n7555 n7567_not ; n7568
g7313 and n7566_not n7567_not ; n7569
g7314 and n7568_not n7569_not ; n7570
g7315 and n7259_not n7261_not ; n7571
g7316 and n7570_not n7571_not ; n7572
g7317 and n7570 n7571 ; n7573
g7318 and n7572_not n7573_not ; n7574
g7319 and n7399_not n7574 ; n7575
g7320 and n7399_not n7575_not ; n7576
g7321 and n7574 n7575_not ; n7577
g7322 and n7576_not n7577_not ; n7578
g7323 and n7388_not n7578_not ; n7579
g7324 and n7388_not n7579_not ; n7580
g7325 and n7578_not n7579_not ; n7581
g7326 and n7580_not n7581_not ; n7582
g7327 and b[31] n1302 ; n7583
g7328 and b[29] n1391 ; n7584
g7329 and b[30] n1297 ; n7585
g7330 and n7584_not n7585_not ; n7586
g7331 and n7583_not n7586 ; n7587
g7332 and n1305 n3796 ; n7588
g7333 and n7587 n7588_not ; n7589
g7334 and a[17] n7589_not ; n7590
g7335 and a[17] n7590_not ; n7591
g7336 and n7589_not n7590_not ; n7592
g7337 and n7591_not n7592_not ; n7593
g7338 and n7582 n7593 ; n7594
g7339 and n7582_not n7593_not ; n7595
g7340 and n7594_not n7595_not ; n7596
g7341 and n7386_not n7596 ; n7597
g7342 and n7386 n7596_not ; n7598
g7343 and n7597_not n7598_not ; n7599
g7344 and n7385_not n7599 ; n7600
g7345 and n7599 n7600_not ; n7601
g7346 and n7385_not n7600_not ; n7602
g7347 and n7601_not n7602_not ; n7603
g7348 and n7088_not n7291_not ; n7604
g7349 and n7288_not n7604_not ; n7605
g7350 and n7603 n7605 ; n7606
g7351 and n7603_not n7605_not ; n7607
g7352 and n7606_not n7607_not ; n7608
g7353 and b[37] n700 ; n7609
g7354 and b[35] n767 ; n7610
g7355 and b[36] n695 ; n7611
g7356 and n7610_not n7611_not ; n7612
g7357 and n7609_not n7612 ; n7613
g7358 and n703 n5181 ; n7614
g7359 and n7613 n7614_not ; n7615
g7360 and a[11] n7615_not ; n7616
g7361 and a[11] n7616_not ; n7617
g7362 and n7615_not n7616_not ; n7618
g7363 and n7617_not n7618_not ; n7619
g7364 and n7608 n7619_not ; n7620
g7365 and n7608 n7620_not ; n7621
g7366 and n7619_not n7620_not ; n7622
g7367 and n7621_not n7622_not ; n7623
g7368 and n7306_not n7310_not ; n7624
g7369 and n7623 n7624 ; n7625
g7370 and n7623_not n7624_not ; n7626
g7371 and n7625_not n7626_not ; n7627
g7372 and b[40] n511 ; n7628
g7373 and b[38] n541 ; n7629
g7374 and b[39] n506 ; n7630
g7375 and n7629_not n7630_not ; n7631
g7376 and n7628_not n7631 ; n7632
g7377 and n514 n5955 ; n7633
g7378 and n7632 n7633_not ; n7634
g7379 and a[8] n7634_not ; n7635
g7380 and a[8] n7635_not ; n7636
g7381 and n7634_not n7635_not ; n7637
g7382 and n7636_not n7637_not ; n7638
g7383 and n7627 n7638_not ; n7639
g7384 and n7627_not n7638 ; n7640
g7385 and n7374_not n7640_not ; n7641
g7386 and n7639_not n7641 ; n7642
g7387 and n7374_not n7642_not ; n7643
g7388 and n7639_not n7642_not ; n7644
g7389 and n7640_not n7644 ; n7645
g7390 and n7643_not n7645_not ; n7646
g7391 and b[43] n362 ; n7647
g7392 and b[41] n403 ; n7648
g7393 and b[42] n357 ; n7649
g7394 and n7648_not n7649_not ; n7650
g7395 and n7647_not n7650 ; n7651
g7396 and n365 n6515 ; n7652
g7397 and n7651 n7652_not ; n7653
g7398 and a[5] n7653_not ; n7654
g7399 and a[5] n7654_not ; n7655
g7400 and n7653_not n7654_not ; n7656
g7401 and n7655_not n7656_not ; n7657
g7402 and n7646_not n7657_not ; n7658
g7403 and n7646_not n7658_not ; n7659
g7404 and n7657_not n7658_not ; n7660
g7405 and n7659_not n7660_not ; n7661
g7406 and n7342_not n7348_not ; n7662
g7407 and n7661 n7662 ; n7663
g7408 and n7661_not n7662_not ; n7664
g7409 and n7663_not n7664_not ; n7665
g7410 and b[46] n266 ; n7666
g7411 and b[44] n284 ; n7667
g7412 and b[45] n261 ; n7668
g7413 and n7667_not n7668_not ; n7669
g7414 and n7666_not n7669 ; n7670
g7415 and n7357_not n7359_not ; n7671
g7416 and b[45]_not b[46]_not ; n7672
g7417 and b[45] b[46] ; n7673
g7418 and n7672_not n7673_not ; n7674
g7419 and n7671_not n7674 ; n7675
g7420 and n7671 n7674_not ; n7676
g7421 and n7675_not n7676_not ; n7677
g7422 and n269 n7677 ; n7678
g7423 and n7670 n7678_not ; n7679
g7424 and a[2] n7679_not ; n7680
g7425 and a[2] n7680_not ; n7681
g7426 and n7679_not n7680_not ; n7682
g7427 and n7681_not n7682_not ; n7683
g7428 and n7665 n7683_not ; n7684
g7429 and n7665 n7684_not ; n7685
g7430 and n7683_not n7684_not ; n7686
g7431 and n7685_not n7686_not ; n7687
g7432 and n7369_not n7371_not ; n7688
g7433 and n7687_not n7688_not ; n7689
g7434 and n7687 n7688 ; n7690
g7435 and n7689_not n7690_not ; f[46]
g7436 and b[47] n266 ; n7692
g7437 and b[45] n284 ; n7693
g7438 and b[46] n261 ; n7694
g7439 and n7693_not n7694_not ; n7695
g7440 and n7692_not n7695 ; n7696
g7441 and n7673_not n7675_not ; n7697
g7442 and b[46]_not b[47]_not ; n7698
g7443 and b[46] b[47] ; n7699
g7444 and n7698_not n7699_not ; n7700
g7445 and n7697_not n7700 ; n7701
g7446 and n7697 n7700_not ; n7702
g7447 and n7701_not n7702_not ; n7703
g7448 and n269 n7703 ; n7704
g7449 and n7696 n7704_not ; n7705
g7450 and a[2] n7705_not ; n7706
g7451 and a[2] n7706_not ; n7707
g7452 and n7705_not n7706_not ; n7708
g7453 and n7707_not n7708_not ; n7709
g7454 and n7658_not n7664_not ; n7710
g7455 and b[35] n951 ; n7711
g7456 and b[33] n1056 ; n7712
g7457 and b[34] n946 ; n7713
g7458 and n7712_not n7713_not ; n7714
g7459 and n7711_not n7714 ; n7715
g7460 and n954 n4696 ; n7716
g7461 and n7715 n7716_not ; n7717
g7462 and a[14] n7717_not ; n7718
g7463 and a[14] n7718_not ; n7719
g7464 and n7717_not n7718_not ; n7720
g7465 and n7719_not n7720_not ; n7721
g7466 and n7595_not n7597_not ; n7722
g7467 and b[32] n1302 ; n7723
g7468 and b[30] n1391 ; n7724
g7469 and b[31] n1297 ; n7725
g7470 and n7724_not n7725_not ; n7726
g7471 and n7723_not n7726 ; n7727
g7472 and n1305 n4013 ; n7728
g7473 and n7727 n7728_not ; n7729
g7474 and a[17] n7729_not ; n7730
g7475 and a[17] n7730_not ; n7731
g7476 and n7729_not n7730_not ; n7732
g7477 and n7731_not n7732_not ; n7733
g7478 and n7575_not n7579_not ; n7734
g7479 and b[29] n1627 ; n7735
g7480 and b[27] n1763 ; n7736
g7481 and b[28] n1622 ; n7737
g7482 and n7736_not n7737_not ; n7738
g7483 and n7735_not n7738 ; n7739
g7484 and n1630 n3383 ; n7740
g7485 and n7739 n7740_not ; n7741
g7486 and a[20] n7741_not ; n7742
g7487 and a[20] n7742_not ; n7743
g7488 and n7741_not n7742_not ; n7744
g7489 and n7743_not n7744_not ; n7745
g7490 and n7567_not n7572_not ; n7746
g7491 and n7548_not n7554_not ; n7747
g7492 and n7509_not n7516_not ; n7748
g7493 and b[17] n3638 ; n7749
g7494 and b[15] n3843 ; n7750
g7495 and b[16] n3633 ; n7751
g7496 and n7750_not n7751_not ; n7752
g7497 and n7749_not n7752 ; n7753
g7498 and n1356 n3641 ; n7754
g7499 and n7753 n7754_not ; n7755
g7500 and a[32] n7755_not ; n7756
g7501 and a[32] n7756_not ; n7757
g7502 and n7755_not n7756_not ; n7758
g7503 and n7757_not n7758_not ; n7759
g7504 and n7504_not n7506_not ; n7760
g7505 and b[14] n4287 ; n7761
g7506 and b[12] n4532 ; n7762
g7507 and b[13] n4282 ; n7763
g7508 and n7762_not n7763_not ; n7764
g7509 and n7761_not n7764 ; n7765
g7510 and n1034 n4290 ; n7766
g7511 and n7765 n7766_not ; n7767
g7512 and a[35] n7767_not ; n7768
g7513 and a[35] n7768_not ; n7769
g7514 and n7767_not n7768_not ; n7770
g7515 and n7769_not n7770_not ; n7771
g7516 and n7465_not n7471_not ; n7772
g7517 and b[8] n5777 ; n7773
g7518 and b[6] n6059 ; n7774
g7519 and b[7] n5772 ; n7775
g7520 and n7774_not n7775_not ; n7776
g7521 and n7773_not n7776 ; n7777
g7522 and n585 n5780 ; n7778
g7523 and n7777 n7778_not ; n7779
g7524 and a[41] n7779_not ; n7780
g7525 and a[41] n7780_not ; n7781
g7526 and n7779_not n7780_not ; n7782
g7527 and n7781_not n7782_not ; n7783
g7528 and n7460_not n7462_not ; n7784
g7529 and b[2] n7446 ; n7785
g7530 and n7152 n7445_not ; n7786
g7531 and n7440 n7786 ; n7787
g7532 and b[0] n7787 ; n7788
g7533 and b[1] n7441 ; n7789
g7534 and n7788_not n7789_not ; n7790
g7535 and n7785_not n7790 ; n7791
g7536 and n296 n7449 ; n7792
g7537 and n7791 n7792_not ; n7793
g7538 and a[47] n7793_not ; n7794
g7539 and a[47] n7794_not ; n7795
g7540 and n7793_not n7794_not ; n7796
g7541 and n7795_not n7796_not ; n7797
g7542 and n7456_not n7797 ; n7798
g7543 and n7456 n7797_not ; n7799
g7544 and n7798_not n7799_not ; n7800
g7545 and b[5] n6595 ; n7801
g7546 and b[3] n6902 ; n7802
g7547 and b[4] n6590 ; n7803
g7548 and n7802_not n7803_not ; n7804
g7549 and n7801_not n7804 ; n7805
g7550 and n394 n6598 ; n7806
g7551 and n7805 n7806_not ; n7807
g7552 and a[44] n7807_not ; n7808
g7553 and a[44] n7808_not ; n7809
g7554 and n7807_not n7808_not ; n7810
g7555 and n7809_not n7810_not ; n7811
g7556 and n7800 n7811_not ; n7812
g7557 and n7800 n7812_not ; n7813
g7558 and n7811_not n7812_not ; n7814
g7559 and n7813_not n7814_not ; n7815
g7560 and n7784_not n7815_not ; n7816
g7561 and n7784 n7815 ; n7817
g7562 and n7816_not n7817_not ; n7818
g7563 and n7783_not n7818 ; n7819
g7564 and n7783_not n7819_not ; n7820
g7565 and n7818 n7819_not ; n7821
g7566 and n7820_not n7821_not ; n7822
g7567 and n7772_not n7822_not ; n7823
g7568 and n7772_not n7823_not ; n7824
g7569 and n7822_not n7823_not ; n7825
g7570 and n7824_not n7825_not ; n7826
g7571 and b[11] n5035 ; n7827
g7572 and b[9] n5277 ; n7828
g7573 and b[10] n5030 ; n7829
g7574 and n7828_not n7829_not ; n7830
g7575 and n7827_not n7830 ; n7831
g7576 and n818 n5038 ; n7832
g7577 and n7831 n7832_not ; n7833
g7578 and a[38] n7833_not ; n7834
g7579 and a[38] n7834_not ; n7835
g7580 and n7833_not n7834_not ; n7836
g7581 and n7835_not n7836_not ; n7837
g7582 and n7826 n7837 ; n7838
g7583 and n7826_not n7837_not ; n7839
g7584 and n7838_not n7839_not ; n7840
g7585 and n7489_not n7840 ; n7841
g7586 and n7489 n7840_not ; n7842
g7587 and n7841_not n7842_not ; n7843
g7588 and n7771_not n7843 ; n7844
g7589 and n7843 n7844_not ; n7845
g7590 and n7771_not n7844_not ; n7846
g7591 and n7845_not n7846_not ; n7847
g7592 and n7760_not n7847_not ; n7848
g7593 and n7760 n7847 ; n7849
g7594 and n7848_not n7849_not ; n7850
g7595 and n7759_not n7850 ; n7851
g7596 and n7759_not n7851_not ; n7852
g7597 and n7850 n7851_not ; n7853
g7598 and n7852_not n7853_not ; n7854
g7599 and n7748_not n7854_not ; n7855
g7600 and n7748_not n7855_not ; n7856
g7601 and n7854_not n7855_not ; n7857
g7602 and n7856_not n7857_not ; n7858
g7603 and b[20] n3050 ; n7859
g7604 and b[18] n3243 ; n7860
g7605 and b[19] n3045 ; n7861
g7606 and n7860_not n7861_not ; n7862
g7607 and n7859_not n7862 ; n7863
g7608 and n1846 n3053 ; n7864
g7609 and n7863 n7864_not ; n7865
g7610 and a[29] n7865_not ; n7866
g7611 and a[29] n7866_not ; n7867
g7612 and n7865_not n7866_not ; n7868
g7613 and n7867_not n7868_not ; n7869
g7614 and n7858_not n7869_not ; n7870
g7615 and n7858_not n7870_not ; n7871
g7616 and n7869_not n7870_not ; n7872
g7617 and n7871_not n7872_not ; n7873
g7618 and n7529_not n7535_not ; n7874
g7619 and n7873 n7874 ; n7875
g7620 and n7873_not n7874_not ; n7876
g7621 and n7875_not n7876_not ; n7877
g7622 and b[23] n2539 ; n7878
g7623 and b[21] n2685 ; n7879
g7624 and b[22] n2534 ; n7880
g7625 and n7879_not n7880_not ; n7881
g7626 and n7878_not n7881 ; n7882
g7627 and n2300 n2542 ; n7883
g7628 and n7882 n7883_not ; n7884
g7629 and a[26] n7884_not ; n7885
g7630 and a[26] n7885_not ; n7886
g7631 and n7884_not n7885_not ; n7887
g7632 and n7886_not n7887_not ; n7888
g7633 and n7877 n7888_not ; n7889
g7634 and n7877_not n7888 ; n7890
g7635 and n7747_not n7890_not ; n7891
g7636 and n7889_not n7891 ; n7892
g7637 and n7747_not n7892_not ; n7893
g7638 and n7889_not n7892_not ; n7894
g7639 and n7890_not n7894 ; n7895
g7640 and n7893_not n7895_not ; n7896
g7641 and b[26] n2048 ; n7897
g7642 and b[24] n2198 ; n7898
g7643 and b[25] n2043 ; n7899
g7644 and n7898_not n7899_not ; n7900
g7645 and n7897_not n7900 ; n7901
g7646 and n2051 n2813 ; n7902
g7647 and n7901 n7902_not ; n7903
g7648 and a[23] n7903_not ; n7904
g7649 and a[23] n7904_not ; n7905
g7650 and n7903_not n7904_not ; n7906
g7651 and n7905_not n7906_not ; n7907
g7652 and n7896 n7907 ; n7908
g7653 and n7896_not n7907_not ; n7909
g7654 and n7908_not n7909_not ; n7910
g7655 and n7746_not n7910 ; n7911
g7656 and n7746 n7910_not ; n7912
g7657 and n7911_not n7912_not ; n7913
g7658 and n7745 n7913_not ; n7914
g7659 and n7745_not n7913 ; n7915
g7660 and n7914_not n7915_not ; n7916
g7661 and n7734_not n7916 ; n7917
g7662 and n7734 n7916_not ; n7918
g7663 and n7917_not n7918_not ; n7919
g7664 and n7733 n7919_not ; n7920
g7665 and n7733_not n7919 ; n7921
g7666 and n7920_not n7921_not ; n7922
g7667 and n7722_not n7922 ; n7923
g7668 and n7722 n7922_not ; n7924
g7669 and n7923_not n7924_not ; n7925
g7670 and n7721_not n7925 ; n7926
g7671 and n7925 n7926_not ; n7927
g7672 and n7721_not n7926_not ; n7928
g7673 and n7927_not n7928_not ; n7929
g7674 and n7600_not n7607_not ; n7930
g7675 and n7929 n7930 ; n7931
g7676 and n7929_not n7930_not ; n7932
g7677 and n7931_not n7932_not ; n7933
g7678 and b[38] n700 ; n7934
g7679 and b[36] n767 ; n7935
g7680 and b[37] n695 ; n7936
g7681 and n7935_not n7936_not ; n7937
g7682 and n7934_not n7937 ; n7938
g7683 and n703 n5205 ; n7939
g7684 and n7938 n7939_not ; n7940
g7685 and a[11] n7940_not ; n7941
g7686 and a[11] n7941_not ; n7942
g7687 and n7940_not n7941_not ; n7943
g7688 and n7942_not n7943_not ; n7944
g7689 and n7933 n7944_not ; n7945
g7690 and n7933 n7945_not ; n7946
g7691 and n7944_not n7945_not ; n7947
g7692 and n7946_not n7947_not ; n7948
g7693 and n7620_not n7626_not ; n7949
g7694 and n7948 n7949 ; n7950
g7695 and n7948_not n7949_not ; n7951
g7696 and n7950_not n7951_not ; n7952
g7697 and b[41] n511 ; n7953
g7698 and b[39] n541 ; n7954
g7699 and b[40] n506 ; n7955
g7700 and n7954_not n7955_not ; n7956
g7701 and n7953_not n7956 ; n7957
g7702 and n514 n6219 ; n7958
g7703 and n7957 n7958_not ; n7959
g7704 and a[8] n7959_not ; n7960
g7705 and a[8] n7960_not ; n7961
g7706 and n7959_not n7960_not ; n7962
g7707 and n7961_not n7962_not ; n7963
g7708 and n7952 n7963_not ; n7964
g7709 and n7952_not n7963 ; n7965
g7710 and n7644_not n7965_not ; n7966
g7711 and n7964_not n7966 ; n7967
g7712 and n7644_not n7967_not ; n7968
g7713 and n7964_not n7967_not ; n7969
g7714 and n7965_not n7969 ; n7970
g7715 and n7968_not n7970_not ; n7971
g7716 and b[44] n362 ; n7972
g7717 and b[42] n403 ; n7973
g7718 and b[43] n357 ; n7974
g7719 and n7973_not n7974_not ; n7975
g7720 and n7972_not n7975 ; n7976
g7721 and n365 n7072 ; n7977
g7722 and n7976 n7977_not ; n7978
g7723 and a[5] n7978_not ; n7979
g7724 and a[5] n7979_not ; n7980
g7725 and n7978_not n7979_not ; n7981
g7726 and n7980_not n7981_not ; n7982
g7727 and n7971 n7982 ; n7983
g7728 and n7971_not n7982_not ; n7984
g7729 and n7983_not n7984_not ; n7985
g7730 and n7710_not n7985 ; n7986
g7731 and n7710 n7985_not ; n7987
g7732 and n7986_not n7987_not ; n7988
g7733 and n7709_not n7988 ; n7989
g7734 and n7988 n7989_not ; n7990
g7735 and n7709_not n7989_not ; n7991
g7736 and n7990_not n7991_not ; n7992
g7737 and n7684_not n7689_not ; n7993
g7738 and n7992_not n7993_not ; n7994
g7739 and n7992 n7993 ; n7995
g7740 and n7994_not n7995_not ; f[47]
g7741 and n7989_not n7994_not ; n7997
g7742 and b[48] n266 ; n7998
g7743 and b[46] n284 ; n7999
g7744 and b[47] n261 ; n8000
g7745 and n7999_not n8000_not ; n8001
g7746 and n7998_not n8001 ; n8002
g7747 and n7699_not n7701_not ; n8003
g7748 and b[47]_not b[48]_not ; n8004
g7749 and b[47] b[48] ; n8005
g7750 and n8004_not n8005_not ; n8006
g7751 and n8003_not n8006 ; n8007
g7752 and n8003 n8006_not ; n8008
g7753 and n8007_not n8008_not ; n8009
g7754 and n269 n8009 ; n8010
g7755 and n8002 n8010_not ; n8011
g7756 and a[2] n8011_not ; n8012
g7757 and a[2] n8012_not ; n8013
g7758 and n8011_not n8012_not ; n8014
g7759 and n8013_not n8014_not ; n8015
g7760 and n7984_not n7986_not ; n8016
g7761 and n7926_not n7932_not ; n8017
g7762 and n7921_not n7923_not ; n8018
g7763 and b[33] n1302 ; n8019
g7764 and b[31] n1391 ; n8020
g7765 and b[32] n1297 ; n8021
g7766 and n8020_not n8021_not ; n8022
g7767 and n8019_not n8022 ; n8023
g7768 and n1305 n4223 ; n8024
g7769 and n8023 n8024_not ; n8025
g7770 and a[17] n8025_not ; n8026
g7771 and a[17] n8026_not ; n8027
g7772 and n8025_not n8026_not ; n8028
g7773 and n8027_not n8028_not ; n8029
g7774 and n7915_not n7917_not ; n8030
g7775 and n7909_not n7911_not ; n8031
g7776 and b[27] n2048 ; n8032
g7777 and b[25] n2198 ; n8033
g7778 and b[26] n2043 ; n8034
g7779 and n8033_not n8034_not ; n8035
g7780 and n8032_not n8035 ; n8036
g7781 and n2051 n2990 ; n8037
g7782 and n8036 n8037_not ; n8038
g7783 and a[23] n8038_not ; n8039
g7784 and a[23] n8039_not ; n8040
g7785 and n8038_not n8039_not ; n8041
g7786 and n8040_not n8041_not ; n8042
g7787 and n7844_not n7848_not ; n8043
g7788 and b[15] n4287 ; n8044
g7789 and b[13] n4532 ; n8045
g7790 and b[14] n4282 ; n8046
g7791 and n8045_not n8046_not ; n8047
g7792 and n8044_not n8047 ; n8048
g7793 and n1131 n4290 ; n8049
g7794 and n8048 n8049_not ; n8050
g7795 and a[35] n8050_not ; n8051
g7796 and a[35] n8051_not ; n8052
g7797 and n8050_not n8051_not ; n8053
g7798 and n8052_not n8053_not ; n8054
g7799 and n7839_not n7841_not ; n8055
g7800 and b[12] n5035 ; n8056
g7801 and b[10] n5277 ; n8057
g7802 and b[11] n5030 ; n8058
g7803 and n8057_not n8058_not ; n8059
g7804 and n8056_not n8059 ; n8060
g7805 and n842 n5038 ; n8061
g7806 and n8060 n8061_not ; n8062
g7807 and a[38] n8062_not ; n8063
g7808 and a[38] n8063_not ; n8064
g7809 and n8062_not n8063_not ; n8065
g7810 and n8064_not n8065_not ; n8066
g7811 and n7819_not n7823_not ; n8067
g7812 and b[6] n6595 ; n8068
g7813 and b[4] n6902 ; n8069
g7814 and b[5] n6590 ; n8070
g7815 and n8069_not n8070_not ; n8071
g7816 and n8068_not n8071 ; n8072
g7817 and n459 n6598 ; n8073
g7818 and n8072 n8073_not ; n8074
g7819 and a[44] n8074_not ; n8075
g7820 and a[44] n8075_not ; n8076
g7821 and n8074_not n8075_not ; n8077
g7822 and n8076_not n8077_not ; n8078
g7823 and a[47] a[48]_not ; n8079
g7824 and a[47]_not a[48] ; n8080
g7825 and n8079_not n8080_not ; n8081
g7826 and b[0] n8081_not ; n8082
g7827 and n7799_not n8082 ; n8083
g7828 and n7799 n8082_not ; n8084
g7829 and n8083_not n8084_not ; n8085
g7830 and b[3] n7446 ; n8086
g7831 and b[1] n7787 ; n8087
g7832 and b[2] n7441 ; n8088
g7833 and n8087_not n8088_not ; n8089
g7834 and n8086_not n8089 ; n8090
g7835 and n318 n7449 ; n8091
g7836 and n8090 n8091_not ; n8092
g7837 and a[47] n8092_not ; n8093
g7838 and a[47] n8093_not ; n8094
g7839 and n8092_not n8093_not ; n8095
g7840 and n8094_not n8095_not ; n8096
g7841 and n8085_not n8096_not ; n8097
g7842 and n8085 n8096 ; n8098
g7843 and n8097_not n8098_not ; n8099
g7844 and n8078_not n8099 ; n8100
g7845 and n8099 n8100_not ; n8101
g7846 and n8078_not n8100_not ; n8102
g7847 and n8101_not n8102_not ; n8103
g7848 and n7812_not n7816_not ; n8104
g7849 and n8103 n8104 ; n8105
g7850 and n8103_not n8104_not ; n8106
g7851 and n8105_not n8106_not ; n8107
g7852 and b[9] n5777 ; n8108
g7853 and b[7] n6059 ; n8109
g7854 and b[8] n5772 ; n8110
g7855 and n8109_not n8110_not ; n8111
g7856 and n8108_not n8111 ; n8112
g7857 and n651 n5780 ; n8113
g7858 and n8112 n8113_not ; n8114
g7859 and a[41] n8114_not ; n8115
g7860 and a[41] n8115_not ; n8116
g7861 and n8114_not n8115_not ; n8117
g7862 and n8116_not n8117_not ; n8118
g7863 and n8107_not n8118 ; n8119
g7864 and n8107 n8118_not ; n8120
g7865 and n8119_not n8120_not ; n8121
g7866 and n8067_not n8121 ; n8122
g7867 and n8067 n8121_not ; n8123
g7868 and n8122_not n8123_not ; n8124
g7869 and n8066_not n8124 ; n8125
g7870 and n8066_not n8125_not ; n8126
g7871 and n8124 n8125_not ; n8127
g7872 and n8126_not n8127_not ; n8128
g7873 and n8055_not n8128_not ; n8129
g7874 and n8055 n8127_not ; n8130
g7875 and n8126_not n8130 ; n8131
g7876 and n8129_not n8131_not ; n8132
g7877 and n8054_not n8132 ; n8133
g7878 and n8054 n8132_not ; n8134
g7879 and n8133_not n8134_not ; n8135
g7880 and n8043_not n8135 ; n8136
g7881 and n8043 n8135_not ; n8137
g7882 and n8136_not n8137_not ; n8138
g7883 and b[18] n3638 ; n8139
g7884 and b[16] n3843 ; n8140
g7885 and b[17] n3633 ; n8141
g7886 and n8140_not n8141_not ; n8142
g7887 and n8139_not n8142 ; n8143
g7888 and n1566 n3641 ; n8144
g7889 and n8143 n8144_not ; n8145
g7890 and a[32] n8145_not ; n8146
g7891 and a[32] n8146_not ; n8147
g7892 and n8145_not n8146_not ; n8148
g7893 and n8147_not n8148_not ; n8149
g7894 and n8138 n8149_not ; n8150
g7895 and n8138 n8150_not ; n8151
g7896 and n8149_not n8150_not ; n8152
g7897 and n8151_not n8152_not ; n8153
g7898 and n7851_not n7855_not ; n8154
g7899 and n8153 n8154 ; n8155
g7900 and n8153_not n8154_not ; n8156
g7901 and n8155_not n8156_not ; n8157
g7902 and b[21] n3050 ; n8158
g7903 and b[19] n3243 ; n8159
g7904 and b[20] n3045 ; n8160
g7905 and n8159_not n8160_not ; n8161
g7906 and n8158_not n8161 ; n8162
g7907 and n1984 n3053 ; n8163
g7908 and n8162 n8163_not ; n8164
g7909 and a[29] n8164_not ; n8165
g7910 and a[29] n8165_not ; n8166
g7911 and n8164_not n8165_not ; n8167
g7912 and n8166_not n8167_not ; n8168
g7913 and n8157 n8168_not ; n8169
g7914 and n8157 n8169_not ; n8170
g7915 and n8168_not n8169_not ; n8171
g7916 and n8170_not n8171_not ; n8172
g7917 and n7870_not n7876_not ; n8173
g7918 and n8172 n8173 ; n8174
g7919 and n8172_not n8173_not ; n8175
g7920 and n8174_not n8175_not ; n8176
g7921 and b[24] n2539 ; n8177
g7922 and b[22] n2685 ; n8178
g7923 and b[23] n2534 ; n8179
g7924 and n8178_not n8179_not ; n8180
g7925 and n8177_not n8180 ; n8181
g7926 and n2458 n2542 ; n8182
g7927 and n8181 n8182_not ; n8183
g7928 and a[26] n8183_not ; n8184
g7929 and a[26] n8184_not ; n8185
g7930 and n8183_not n8184_not ; n8186
g7931 and n8185_not n8186_not ; n8187
g7932 and n8176_not n8187 ; n8188
g7933 and n8176 n8187_not ; n8189
g7934 and n8188_not n8189_not ; n8190
g7935 and n7894_not n8190 ; n8191
g7936 and n7894 n8190_not ; n8192
g7937 and n8191_not n8192_not ; n8193
g7938 and n8042_not n8193 ; n8194
g7939 and n8193 n8194_not ; n8195
g7940 and n8042_not n8194_not ; n8196
g7941 and n8195_not n8196_not ; n8197
g7942 and n8031_not n8197 ; n8198
g7943 and n8031 n8197_not ; n8199
g7944 and n8198_not n8199_not ; n8200
g7945 and b[30] n1627 ; n8201
g7946 and b[28] n1763 ; n8202
g7947 and b[29] n1622 ; n8203
g7948 and n8202_not n8203_not ; n8204
g7949 and n8201_not n8204 ; n8205
g7950 and n1630 n3577 ; n8206
g7951 and n8205 n8206_not ; n8207
g7952 and a[20] n8207_not ; n8208
g7953 and a[20] n8208_not ; n8209
g7954 and n8207_not n8208_not ; n8210
g7955 and n8209_not n8210_not ; n8211
g7956 and n8200_not n8211_not ; n8212
g7957 and n8200 n8211 ; n8213
g7958 and n8212_not n8213_not ; n8214
g7959 and n8030_not n8214 ; n8215
g7960 and n8030 n8214_not ; n8216
g7961 and n8215_not n8216_not ; n8217
g7962 and n8029_not n8217 ; n8218
g7963 and n8217 n8218_not ; n8219
g7964 and n8029_not n8218_not ; n8220
g7965 and n8219_not n8220_not ; n8221
g7966 and n8018_not n8221 ; n8222
g7967 and n8018 n8221_not ; n8223
g7968 and n8222_not n8223_not ; n8224
g7969 and b[36] n951 ; n8225
g7970 and b[34] n1056 ; n8226
g7971 and b[35] n946 ; n8227
g7972 and n8226_not n8227_not ; n8228
g7973 and n8225_not n8228 ; n8229
g7974 and n954 n4922 ; n8230
g7975 and n8229 n8230_not ; n8231
g7976 and a[14] n8231_not ; n8232
g7977 and a[14] n8232_not ; n8233
g7978 and n8231_not n8232_not ; n8234
g7979 and n8233_not n8234_not ; n8235
g7980 and n8224_not n8235_not ; n8236
g7981 and n8224 n8235 ; n8237
g7982 and n8236_not n8237_not ; n8238
g7983 and n8017 n8238_not ; n8239
g7984 and n8017_not n8238 ; n8240
g7985 and n8239_not n8240_not ; n8241
g7986 and b[39] n700 ; n8242
g7987 and b[37] n767 ; n8243
g7988 and b[38] n695 ; n8244
g7989 and n8243_not n8244_not ; n8245
g7990 and n8242_not n8245 ; n8246
g7991 and n703 n5451 ; n8247
g7992 and n8246 n8247_not ; n8248
g7993 and a[11] n8248_not ; n8249
g7994 and a[11] n8249_not ; n8250
g7995 and n8248_not n8249_not ; n8251
g7996 and n8250_not n8251_not ; n8252
g7997 and n8241 n8252_not ; n8253
g7998 and n8241 n8253_not ; n8254
g7999 and n8252_not n8253_not ; n8255
g8000 and n8254_not n8255_not ; n8256
g8001 and n7945_not n7951_not ; n8257
g8002 and n8256 n8257 ; n8258
g8003 and n8256_not n8257_not ; n8259
g8004 and n8258_not n8259_not ; n8260
g8005 and b[42] n511 ; n8261
g8006 and b[40] n541 ; n8262
g8007 and b[41] n506 ; n8263
g8008 and n8262_not n8263_not ; n8264
g8009 and n8261_not n8264 ; n8265
g8010 and n514 n6489 ; n8266
g8011 and n8265 n8266_not ; n8267
g8012 and a[8] n8267_not ; n8268
g8013 and a[8] n8268_not ; n8269
g8014 and n8267_not n8268_not ; n8270
g8015 and n8269_not n8270_not ; n8271
g8016 and n8260 n8271_not ; n8272
g8017 and n8260 n8272_not ; n8273
g8018 and n8271_not n8272_not ; n8274
g8019 and n8273_not n8274_not ; n8275
g8020 and n7969_not n8275 ; n8276
g8021 and n7969 n8275_not ; n8277
g8022 and n8276_not n8277_not ; n8278
g8023 and b[45] n362 ; n8279
g8024 and b[43] n403 ; n8280
g8025 and b[44] n357 ; n8281
g8026 and n8280_not n8281_not ; n8282
g8027 and n8279_not n8282 ; n8283
g8028 and n365 n7361 ; n8284
g8029 and n8283 n8284_not ; n8285
g8030 and a[5] n8285_not ; n8286
g8031 and a[5] n8286_not ; n8287
g8032 and n8285_not n8286_not ; n8288
g8033 and n8287_not n8288_not ; n8289
g8034 and n8278_not n8289_not ; n8290
g8035 and n8278 n8289 ; n8291
g8036 and n8290_not n8291_not ; n8292
g8037 and n8016_not n8292 ; n8293
g8038 and n8016 n8292_not ; n8294
g8039 and n8293_not n8294_not ; n8295
g8040 and n8015 n8295_not ; n8296
g8041 and n8015_not n8295 ; n8297
g8042 and n8296_not n8297_not ; n8298
g8043 and n7997_not n8298 ; n8299
g8044 and n7997 n8298_not ; n8300
g8045 and n8299_not n8300_not ; f[48]
g8046 and n8297_not n8299_not ; n8302
g8047 and n8031_not n8197_not ; n8303
g8048 and n8194_not n8303_not ; n8304
g8049 and b[28] n2048 ; n8305
g8050 and b[26] n2198 ; n8306
g8051 and b[27] n2043 ; n8307
g8052 and n8306_not n8307_not ; n8308
g8053 and n8305_not n8308 ; n8309
g8054 and n2051 n3189 ; n8310
g8055 and n8309 n8310_not ; n8311
g8056 and a[23] n8311_not ; n8312
g8057 and a[23] n8312_not ; n8313
g8058 and n8311_not n8312_not ; n8314
g8059 and n8313_not n8314_not ; n8315
g8060 and b[16] n4287 ; n8316
g8061 and b[14] n4532 ; n8317
g8062 and b[15] n4282 ; n8318
g8063 and n8317_not n8318_not ; n8319
g8064 and n8316_not n8319 ; n8320
g8065 and n1237 n4290 ; n8321
g8066 and n8320 n8321_not ; n8322
g8067 and a[35] n8322_not ; n8323
g8068 and a[35] n8323_not ; n8324
g8069 and n8322_not n8323_not ; n8325
g8070 and n8324_not n8325_not ; n8326
g8071 and n8125_not n8129_not ; n8327
g8072 and n8120_not n8122_not ; n8328
g8073 and b[7] n6595 ; n8329
g8074 and b[5] n6902 ; n8330
g8075 and b[6] n6590 ; n8331
g8076 and n8330_not n8331_not ; n8332
g8077 and n8329_not n8332 ; n8333
g8078 and n484 n6598 ; n8334
g8079 and n8333 n8334_not ; n8335
g8080 and a[44] n8335_not ; n8336
g8081 and a[44] n8336_not ; n8337
g8082 and n8335_not n8336_not ; n8338
g8083 and n8337_not n8338_not ; n8339
g8084 and n7799 n8082 ; n8340
g8085 and n8097_not n8340_not ; n8341
g8086 and b[4] n7446 ; n8342
g8087 and b[2] n7787 ; n8343
g8088 and b[3] n7441 ; n8344
g8089 and n8343_not n8344_not ; n8345
g8090 and n8342_not n8345 ; n8346
g8091 and n346 n7449 ; n8347
g8092 and n8346 n8347_not ; n8348
g8093 and a[47] n8348_not ; n8349
g8094 and a[47] n8349_not ; n8350
g8095 and n8348_not n8349_not ; n8351
g8096 and n8350_not n8351_not ; n8352
g8097 and a[50] n8082_not ; n8353
g8098 and a[48]_not a[49] ; n8354
g8099 and a[48] a[49]_not ; n8355
g8100 and n8354_not n8355_not ; n8356
g8101 and n8081 n8356_not ; n8357
g8102 and b[0] n8357 ; n8358
g8103 and a[49]_not a[50] ; n8359
g8104 and a[49] a[50]_not ; n8360
g8105 and n8359_not n8360_not ; n8361
g8106 and n8081_not n8361 ; n8362
g8107 and b[1] n8362 ; n8363
g8108 and n8358_not n8363_not ; n8364
g8109 and n8081_not n8361_not ; n8365
g8110 and n272_not n8365 ; n8366
g8111 and n8364 n8366_not ; n8367
g8112 and a[50] n8367_not ; n8368
g8113 and a[50] n8368_not ; n8369
g8114 and n8367_not n8368_not ; n8370
g8115 and n8369_not n8370_not ; n8371
g8116 and n8353 n8371_not ; n8372
g8117 and n8353_not n8371 ; n8373
g8118 and n8372_not n8373_not ; n8374
g8119 and n8352 n8374_not ; n8375
g8120 and n8352_not n8374 ; n8376
g8121 and n8375_not n8376_not ; n8377
g8122 and n8341_not n8377 ; n8378
g8123 and n8341 n8377_not ; n8379
g8124 and n8378_not n8379_not ; n8380
g8125 and n8339_not n8380 ; n8381
g8126 and n8380 n8381_not ; n8382
g8127 and n8339_not n8381_not ; n8383
g8128 and n8382_not n8383_not ; n8384
g8129 and n8100_not n8106_not ; n8385
g8130 and n8384 n8385 ; n8386
g8131 and n8384_not n8385_not ; n8387
g8132 and n8386_not n8387_not ; n8388
g8133 and b[10] n5777 ; n8389
g8134 and b[8] n6059 ; n8390
g8135 and b[9] n5772 ; n8391
g8136 and n8390_not n8391_not ; n8392
g8137 and n8389_not n8392 ; n8393
g8138 and n738 n5780 ; n8394
g8139 and n8393 n8394_not ; n8395
g8140 and a[41] n8395_not ; n8396
g8141 and a[41] n8396_not ; n8397
g8142 and n8395_not n8396_not ; n8398
g8143 and n8397_not n8398_not ; n8399
g8144 and n8388 n8399_not ; n8400
g8145 and n8388_not n8399 ; n8401
g8146 and n8328_not n8401_not ; n8402
g8147 and n8400_not n8402 ; n8403
g8148 and n8328_not n8403_not ; n8404
g8149 and n8400_not n8403_not ; n8405
g8150 and n8401_not n8405 ; n8406
g8151 and n8404_not n8406_not ; n8407
g8152 and b[13] n5035 ; n8408
g8153 and b[11] n5277 ; n8409
g8154 and b[12] n5030 ; n8410
g8155 and n8409_not n8410_not ; n8411
g8156 and n8408_not n8411 ; n8412
g8157 and n1008 n5038 ; n8413
g8158 and n8412 n8413_not ; n8414
g8159 and a[38] n8414_not ; n8415
g8160 and a[38] n8415_not ; n8416
g8161 and n8414_not n8415_not ; n8417
g8162 and n8416_not n8417_not ; n8418
g8163 and n8407 n8418 ; n8419
g8164 and n8407_not n8418_not ; n8420
g8165 and n8419_not n8420_not ; n8421
g8166 and n8327_not n8421 ; n8422
g8167 and n8327 n8421_not ; n8423
g8168 and n8422_not n8423_not ; n8424
g8169 and n8326_not n8424 ; n8425
g8170 and n8424 n8425_not ; n8426
g8171 and n8326_not n8425_not ; n8427
g8172 and n8426_not n8427_not ; n8428
g8173 and n8133_not n8136_not ; n8429
g8174 and n8428 n8429 ; n8430
g8175 and n8428_not n8429_not ; n8431
g8176 and n8430_not n8431_not ; n8432
g8177 and b[19] n3638 ; n8433
g8178 and b[17] n3843 ; n8434
g8179 and b[18] n3633 ; n8435
g8180 and n8434_not n8435_not ; n8436
g8181 and n8433_not n8436 ; n8437
g8182 and n1708 n3641 ; n8438
g8183 and n8437 n8438_not ; n8439
g8184 and a[32] n8439_not ; n8440
g8185 and a[32] n8440_not ; n8441
g8186 and n8439_not n8440_not ; n8442
g8187 and n8441_not n8442_not ; n8443
g8188 and n8432 n8443_not ; n8444
g8189 and n8432 n8444_not ; n8445
g8190 and n8443_not n8444_not ; n8446
g8191 and n8445_not n8446_not ; n8447
g8192 and n8150_not n8156_not ; n8448
g8193 and n8447 n8448 ; n8449
g8194 and n8447_not n8448_not ; n8450
g8195 and n8449_not n8450_not ; n8451
g8196 and b[22] n3050 ; n8452
g8197 and b[20] n3243 ; n8453
g8198 and b[21] n3045 ; n8454
g8199 and n8453_not n8454_not ; n8455
g8200 and n8452_not n8455 ; n8456
g8201 and n2145 n3053 ; n8457
g8202 and n8456 n8457_not ; n8458
g8203 and a[29] n8458_not ; n8459
g8204 and a[29] n8459_not ; n8460
g8205 and n8458_not n8459_not ; n8461
g8206 and n8460_not n8461_not ; n8462
g8207 and n8451 n8462_not ; n8463
g8208 and n8451 n8463_not ; n8464
g8209 and n8462_not n8463_not ; n8465
g8210 and n8464_not n8465_not ; n8466
g8211 and n8169_not n8175_not ; n8467
g8212 and n8466 n8467 ; n8468
g8213 and n8466_not n8467_not ; n8469
g8214 and n8468_not n8469_not ; n8470
g8215 and b[25] n2539 ; n8471
g8216 and b[23] n2685 ; n8472
g8217 and b[24] n2534 ; n8473
g8218 and n8472_not n8473_not ; n8474
g8219 and n8471_not n8474 ; n8475
g8220 and n2485 n2542 ; n8476
g8221 and n8475 n8476_not ; n8477
g8222 and a[26] n8477_not ; n8478
g8223 and a[26] n8478_not ; n8479
g8224 and n8477_not n8478_not ; n8480
g8225 and n8479_not n8480_not ; n8481
g8226 and n8470 n8481_not ; n8482
g8227 and n8470 n8482_not ; n8483
g8228 and n8481_not n8482_not ; n8484
g8229 and n8483_not n8484_not ; n8485
g8230 and n8189_not n8191_not ; n8486
g8231 and n8485_not n8486_not ; n8487
g8232 and n8485 n8486 ; n8488
g8233 and n8487_not n8488_not ; n8489
g8234 and n8315_not n8489 ; n8490
g8235 and n8315_not n8490_not ; n8491
g8236 and n8489 n8490_not ; n8492
g8237 and n8491_not n8492_not ; n8493
g8238 and n8304_not n8493_not ; n8494
g8239 and n8304_not n8494_not ; n8495
g8240 and n8493_not n8494_not ; n8496
g8241 and n8495_not n8496_not ; n8497
g8242 and b[31] n1627 ; n8498
g8243 and b[29] n1763 ; n8499
g8244 and b[30] n1622 ; n8500
g8245 and n8499_not n8500_not ; n8501
g8246 and n8498_not n8501 ; n8502
g8247 and n1630 n3796 ; n8503
g8248 and n8502 n8503_not ; n8504
g8249 and a[20] n8504_not ; n8505
g8250 and a[20] n8505_not ; n8506
g8251 and n8504_not n8505_not ; n8507
g8252 and n8506_not n8507_not ; n8508
g8253 and n8497_not n8508_not ; n8509
g8254 and n8497_not n8509_not ; n8510
g8255 and n8508_not n8509_not ; n8511
g8256 and n8510_not n8511_not ; n8512
g8257 and n8212_not n8215_not ; n8513
g8258 and n8512 n8513 ; n8514
g8259 and n8512_not n8513_not ; n8515
g8260 and n8514_not n8515_not ; n8516
g8261 and b[34] n1302 ; n8517
g8262 and b[32] n1391 ; n8518
g8263 and b[33] n1297 ; n8519
g8264 and n8518_not n8519_not ; n8520
g8265 and n8517_not n8520 ; n8521
g8266 and n1305 n4466 ; n8522
g8267 and n8521 n8522_not ; n8523
g8268 and a[17] n8523_not ; n8524
g8269 and a[17] n8524_not ; n8525
g8270 and n8523_not n8524_not ; n8526
g8271 and n8525_not n8526_not ; n8527
g8272 and n8516 n8527_not ; n8528
g8273 and n8516 n8528_not ; n8529
g8274 and n8527_not n8528_not ; n8530
g8275 and n8529_not n8530_not ; n8531
g8276 and n8018_not n8221_not ; n8532
g8277 and n8218_not n8532_not ; n8533
g8278 and n8531 n8533 ; n8534
g8279 and n8531_not n8533_not ; n8535
g8280 and n8534_not n8535_not ; n8536
g8281 and b[37] n951 ; n8537
g8282 and b[35] n1056 ; n8538
g8283 and b[36] n946 ; n8539
g8284 and n8538_not n8539_not ; n8540
g8285 and n8537_not n8540 ; n8541
g8286 and n954 n5181 ; n8542
g8287 and n8541 n8542_not ; n8543
g8288 and a[14] n8543_not ; n8544
g8289 and a[14] n8544_not ; n8545
g8290 and n8543_not n8544_not ; n8546
g8291 and n8545_not n8546_not ; n8547
g8292 and n8536 n8547_not ; n8548
g8293 and n8536 n8548_not ; n8549
g8294 and n8547_not n8548_not ; n8550
g8295 and n8549_not n8550_not ; n8551
g8296 and n8236_not n8240_not ; n8552
g8297 and n8551 n8552 ; n8553
g8298 and n8551_not n8552_not ; n8554
g8299 and n8553_not n8554_not ; n8555
g8300 and b[40] n700 ; n8556
g8301 and b[38] n767 ; n8557
g8302 and b[39] n695 ; n8558
g8303 and n8557_not n8558_not ; n8559
g8304 and n8556_not n8559 ; n8560
g8305 and n703 n5955 ; n8561
g8306 and n8560 n8561_not ; n8562
g8307 and a[11] n8562_not ; n8563
g8308 and a[11] n8563_not ; n8564
g8309 and n8562_not n8563_not ; n8565
g8310 and n8564_not n8565_not ; n8566
g8311 and n8555 n8566_not ; n8567
g8312 and n8555 n8567_not ; n8568
g8313 and n8566_not n8567_not ; n8569
g8314 and n8568_not n8569_not ; n8570
g8315 and n8253_not n8259_not ; n8571
g8316 and n8570 n8571 ; n8572
g8317 and n8570_not n8571_not ; n8573
g8318 and n8572_not n8573_not ; n8574
g8319 and b[43] n511 ; n8575
g8320 and b[41] n541 ; n8576
g8321 and b[42] n506 ; n8577
g8322 and n8576_not n8577_not ; n8578
g8323 and n8575_not n8578 ; n8579
g8324 and n514 n6515 ; n8580
g8325 and n8579 n8580_not ; n8581
g8326 and a[8] n8581_not ; n8582
g8327 and a[8] n8582_not ; n8583
g8328 and n8581_not n8582_not ; n8584
g8329 and n8583_not n8584_not ; n8585
g8330 and n8574 n8585_not ; n8586
g8331 and n8574 n8586_not ; n8587
g8332 and n8585_not n8586_not ; n8588
g8333 and n8587_not n8588_not ; n8589
g8334 and n7969_not n8275_not ; n8590
g8335 and n8272_not n8590_not ; n8591
g8336 and n8589 n8591 ; n8592
g8337 and n8589_not n8591_not ; n8593
g8338 and n8592_not n8593_not ; n8594
g8339 and b[46] n362 ; n8595
g8340 and b[44] n403 ; n8596
g8341 and b[45] n357 ; n8597
g8342 and n8596_not n8597_not ; n8598
g8343 and n8595_not n8598 ; n8599
g8344 and n365 n7677 ; n8600
g8345 and n8599 n8600_not ; n8601
g8346 and a[5] n8601_not ; n8602
g8347 and a[5] n8602_not ; n8603
g8348 and n8601_not n8602_not ; n8604
g8349 and n8603_not n8604_not ; n8605
g8350 and n8594 n8605_not ; n8606
g8351 and n8594 n8606_not ; n8607
g8352 and n8605_not n8606_not ; n8608
g8353 and n8607_not n8608_not ; n8609
g8354 and n8290_not n8293_not ; n8610
g8355 and n8609 n8610 ; n8611
g8356 and n8609_not n8610_not ; n8612
g8357 and n8611_not n8612_not ; n8613
g8358 and b[49] n266 ; n8614
g8359 and b[47] n284 ; n8615
g8360 and b[48] n261 ; n8616
g8361 and n8615_not n8616_not ; n8617
g8362 and n8614_not n8617 ; n8618
g8363 and n8005_not n8007_not ; n8619
g8364 and b[48]_not b[49]_not ; n8620
g8365 and b[48] b[49] ; n8621
g8366 and n8620_not n8621_not ; n8622
g8367 and n8619_not n8622 ; n8623
g8368 and n8619 n8622_not ; n8624
g8369 and n8623_not n8624_not ; n8625
g8370 and n269 n8625 ; n8626
g8371 and n8618 n8626_not ; n8627
g8372 and a[2] n8627_not ; n8628
g8373 and a[2] n8628_not ; n8629
g8374 and n8627_not n8628_not ; n8630
g8375 and n8629_not n8630_not ; n8631
g8376 and n8613_not n8631 ; n8632
g8377 and n8613 n8631_not ; n8633
g8378 and n8632_not n8633_not ; n8634
g8379 and n8302_not n8634 ; n8635
g8380 and n8302 n8634_not ; n8636
g8381 and n8635_not n8636_not ; f[49]
g8382 and n8586_not n8593_not ; n8638
g8383 and b[35] n1302 ; n8639
g8384 and b[33] n1391 ; n8640
g8385 and b[34] n1297 ; n8641
g8386 and n8640_not n8641_not ; n8642
g8387 and n8639_not n8642 ; n8643
g8388 and n1305 n4696 ; n8644
g8389 and n8643 n8644_not ; n8645
g8390 and a[17] n8645_not ; n8646
g8391 and a[17] n8646_not ; n8647
g8392 and n8645_not n8646_not ; n8648
g8393 and n8647_not n8648_not ; n8649
g8394 and n8509_not n8515_not ; n8650
g8395 and b[32] n1627 ; n8651
g8396 and b[30] n1763 ; n8652
g8397 and b[31] n1622 ; n8653
g8398 and n8652_not n8653_not ; n8654
g8399 and n8651_not n8654 ; n8655
g8400 and n1630 n4013 ; n8656
g8401 and n8655 n8656_not ; n8657
g8402 and a[20] n8657_not ; n8658
g8403 and a[20] n8658_not ; n8659
g8404 and n8657_not n8658_not ; n8660
g8405 and n8659_not n8660_not ; n8661
g8406 and n8490_not n8494_not ; n8662
g8407 and b[29] n2048 ; n8663
g8408 and b[27] n2198 ; n8664
g8409 and b[28] n2043 ; n8665
g8410 and n8664_not n8665_not ; n8666
g8411 and n8663_not n8666 ; n8667
g8412 and n2051 n3383 ; n8668
g8413 and n8667 n8668_not ; n8669
g8414 and a[23] n8669_not ; n8670
g8415 and a[23] n8670_not ; n8671
g8416 and n8669_not n8670_not ; n8672
g8417 and n8671_not n8672_not ; n8673
g8418 and n8482_not n8487_not ; n8674
g8419 and n8463_not n8469_not ; n8675
g8420 and n8425_not n8431_not ; n8676
g8421 and b[17] n4287 ; n8677
g8422 and b[15] n4532 ; n8678
g8423 and b[16] n4282 ; n8679
g8424 and n8678_not n8679_not ; n8680
g8425 and n8677_not n8680 ; n8681
g8426 and n1356 n4290 ; n8682
g8427 and n8681 n8682_not ; n8683
g8428 and a[35] n8683_not ; n8684
g8429 and a[35] n8684_not ; n8685
g8430 and n8683_not n8684_not ; n8686
g8431 and n8685_not n8686_not ; n8687
g8432 and n8420_not n8422_not ; n8688
g8433 and b[14] n5035 ; n8689
g8434 and b[12] n5277 ; n8690
g8435 and b[13] n5030 ; n8691
g8436 and n8690_not n8691_not ; n8692
g8437 and n8689_not n8692 ; n8693
g8438 and n1034 n5038 ; n8694
g8439 and n8693 n8694_not ; n8695
g8440 and a[38] n8695_not ; n8696
g8441 and a[38] n8696_not ; n8697
g8442 and n8695_not n8696_not ; n8698
g8443 and n8697_not n8698_not ; n8699
g8444 and n8381_not n8387_not ; n8700
g8445 and b[8] n6595 ; n8701
g8446 and b[6] n6902 ; n8702
g8447 and b[7] n6590 ; n8703
g8448 and n8702_not n8703_not ; n8704
g8449 and n8701_not n8704 ; n8705
g8450 and n585 n6598 ; n8706
g8451 and n8705 n8706_not ; n8707
g8452 and a[44] n8707_not ; n8708
g8453 and a[44] n8708_not ; n8709
g8454 and n8707_not n8708_not ; n8710
g8455 and n8709_not n8710_not ; n8711
g8456 and n8376_not n8378_not ; n8712
g8457 and b[2] n8362 ; n8713
g8458 and n8081 n8361_not ; n8714
g8459 and n8356 n8714 ; n8715
g8460 and b[0] n8715 ; n8716
g8461 and b[1] n8357 ; n8717
g8462 and n8716_not n8717_not ; n8718
g8463 and n8713_not n8718 ; n8719
g8464 and n296 n8365 ; n8720
g8465 and n8719 n8720_not ; n8721
g8466 and a[50] n8721_not ; n8722
g8467 and a[50] n8722_not ; n8723
g8468 and n8721_not n8722_not ; n8724
g8469 and n8723_not n8724_not ; n8725
g8470 and n8372_not n8725 ; n8726
g8471 and n8372 n8725_not ; n8727
g8472 and n8726_not n8727_not ; n8728
g8473 and b[5] n7446 ; n8729
g8474 and b[3] n7787 ; n8730
g8475 and b[4] n7441 ; n8731
g8476 and n8730_not n8731_not ; n8732
g8477 and n8729_not n8732 ; n8733
g8478 and n394 n7449 ; n8734
g8479 and n8733 n8734_not ; n8735
g8480 and a[47] n8735_not ; n8736
g8481 and a[47] n8736_not ; n8737
g8482 and n8735_not n8736_not ; n8738
g8483 and n8737_not n8738_not ; n8739
g8484 and n8728 n8739_not ; n8740
g8485 and n8728 n8740_not ; n8741
g8486 and n8739_not n8740_not ; n8742
g8487 and n8741_not n8742_not ; n8743
g8488 and n8712_not n8743_not ; n8744
g8489 and n8712 n8743 ; n8745
g8490 and n8744_not n8745_not ; n8746
g8491 and n8711_not n8746 ; n8747
g8492 and n8711_not n8747_not ; n8748
g8493 and n8746 n8747_not ; n8749
g8494 and n8748_not n8749_not ; n8750
g8495 and n8700_not n8750_not ; n8751
g8496 and n8700_not n8751_not ; n8752
g8497 and n8750_not n8751_not ; n8753
g8498 and n8752_not n8753_not ; n8754
g8499 and b[11] n5777 ; n8755
g8500 and b[9] n6059 ; n8756
g8501 and b[10] n5772 ; n8757
g8502 and n8756_not n8757_not ; n8758
g8503 and n8755_not n8758 ; n8759
g8504 and n818 n5780 ; n8760
g8505 and n8759 n8760_not ; n8761
g8506 and a[41] n8761_not ; n8762
g8507 and a[41] n8762_not ; n8763
g8508 and n8761_not n8762_not ; n8764
g8509 and n8763_not n8764_not ; n8765
g8510 and n8754 n8765 ; n8766
g8511 and n8754_not n8765_not ; n8767
g8512 and n8766_not n8767_not ; n8768
g8513 and n8405_not n8768 ; n8769
g8514 and n8405 n8768_not ; n8770
g8515 and n8769_not n8770_not ; n8771
g8516 and n8699_not n8771 ; n8772
g8517 and n8771 n8772_not ; n8773
g8518 and n8699_not n8772_not ; n8774
g8519 and n8773_not n8774_not ; n8775
g8520 and n8688_not n8775_not ; n8776
g8521 and n8688 n8775 ; n8777
g8522 and n8776_not n8777_not ; n8778
g8523 and n8687_not n8778 ; n8779
g8524 and n8687_not n8779_not ; n8780
g8525 and n8778 n8779_not ; n8781
g8526 and n8780_not n8781_not ; n8782
g8527 and n8676_not n8782_not ; n8783
g8528 and n8676_not n8783_not ; n8784
g8529 and n8782_not n8783_not ; n8785
g8530 and n8784_not n8785_not ; n8786
g8531 and b[20] n3638 ; n8787
g8532 and b[18] n3843 ; n8788
g8533 and b[19] n3633 ; n8789
g8534 and n8788_not n8789_not ; n8790
g8535 and n8787_not n8790 ; n8791
g8536 and n1846 n3641 ; n8792
g8537 and n8791 n8792_not ; n8793
g8538 and a[32] n8793_not ; n8794
g8539 and a[32] n8794_not ; n8795
g8540 and n8793_not n8794_not ; n8796
g8541 and n8795_not n8796_not ; n8797
g8542 and n8786_not n8797_not ; n8798
g8543 and n8786_not n8798_not ; n8799
g8544 and n8797_not n8798_not ; n8800
g8545 and n8799_not n8800_not ; n8801
g8546 and n8444_not n8450_not ; n8802
g8547 and n8801 n8802 ; n8803
g8548 and n8801_not n8802_not ; n8804
g8549 and n8803_not n8804_not ; n8805
g8550 and b[23] n3050 ; n8806
g8551 and b[21] n3243 ; n8807
g8552 and b[22] n3045 ; n8808
g8553 and n8807_not n8808_not ; n8809
g8554 and n8806_not n8809 ; n8810
g8555 and n2300 n3053 ; n8811
g8556 and n8810 n8811_not ; n8812
g8557 and a[29] n8812_not ; n8813
g8558 and a[29] n8813_not ; n8814
g8559 and n8812_not n8813_not ; n8815
g8560 and n8814_not n8815_not ; n8816
g8561 and n8805 n8816_not ; n8817
g8562 and n8805_not n8816 ; n8818
g8563 and n8675_not n8818_not ; n8819
g8564 and n8817_not n8819 ; n8820
g8565 and n8675_not n8820_not ; n8821
g8566 and n8817_not n8820_not ; n8822
g8567 and n8818_not n8822 ; n8823
g8568 and n8821_not n8823_not ; n8824
g8569 and b[26] n2539 ; n8825
g8570 and b[24] n2685 ; n8826
g8571 and b[25] n2534 ; n8827
g8572 and n8826_not n8827_not ; n8828
g8573 and n8825_not n8828 ; n8829
g8574 and n2542 n2813 ; n8830
g8575 and n8829 n8830_not ; n8831
g8576 and a[26] n8831_not ; n8832
g8577 and a[26] n8832_not ; n8833
g8578 and n8831_not n8832_not ; n8834
g8579 and n8833_not n8834_not ; n8835
g8580 and n8824 n8835 ; n8836
g8581 and n8824_not n8835_not ; n8837
g8582 and n8836_not n8837_not ; n8838
g8583 and n8674_not n8838 ; n8839
g8584 and n8674 n8838_not ; n8840
g8585 and n8839_not n8840_not ; n8841
g8586 and n8673 n8841_not ; n8842
g8587 and n8673_not n8841 ; n8843
g8588 and n8842_not n8843_not ; n8844
g8589 and n8662_not n8844 ; n8845
g8590 and n8662 n8844_not ; n8846
g8591 and n8845_not n8846_not ; n8847
g8592 and n8661 n8847_not ; n8848
g8593 and n8661_not n8847 ; n8849
g8594 and n8848_not n8849_not ; n8850
g8595 and n8650_not n8850 ; n8851
g8596 and n8650 n8850_not ; n8852
g8597 and n8851_not n8852_not ; n8853
g8598 and n8649_not n8853 ; n8854
g8599 and n8853 n8854_not ; n8855
g8600 and n8649_not n8854_not ; n8856
g8601 and n8855_not n8856_not ; n8857
g8602 and n8528_not n8535_not ; n8858
g8603 and n8857 n8858 ; n8859
g8604 and n8857_not n8858_not ; n8860
g8605 and n8859_not n8860_not ; n8861
g8606 and b[38] n951 ; n8862
g8607 and b[36] n1056 ; n8863
g8608 and b[37] n946 ; n8864
g8609 and n8863_not n8864_not ; n8865
g8610 and n8862_not n8865 ; n8866
g8611 and n954 n5205 ; n8867
g8612 and n8866 n8867_not ; n8868
g8613 and a[14] n8868_not ; n8869
g8614 and a[14] n8869_not ; n8870
g8615 and n8868_not n8869_not ; n8871
g8616 and n8870_not n8871_not ; n8872
g8617 and n8861 n8872_not ; n8873
g8618 and n8861 n8873_not ; n8874
g8619 and n8872_not n8873_not ; n8875
g8620 and n8874_not n8875_not ; n8876
g8621 and n8548_not n8554_not ; n8877
g8622 and n8876 n8877 ; n8878
g8623 and n8876_not n8877_not ; n8879
g8624 and n8878_not n8879_not ; n8880
g8625 and b[41] n700 ; n8881
g8626 and b[39] n767 ; n8882
g8627 and b[40] n695 ; n8883
g8628 and n8882_not n8883_not ; n8884
g8629 and n8881_not n8884 ; n8885
g8630 and n703 n6219 ; n8886
g8631 and n8885 n8886_not ; n8887
g8632 and a[11] n8887_not ; n8888
g8633 and a[11] n8888_not ; n8889
g8634 and n8887_not n8888_not ; n8890
g8635 and n8889_not n8890_not ; n8891
g8636 and n8880 n8891_not ; n8892
g8637 and n8880 n8892_not ; n8893
g8638 and n8891_not n8892_not ; n8894
g8639 and n8893_not n8894_not ; n8895
g8640 and n8567_not n8573_not ; n8896
g8641 and n8895 n8896 ; n8897
g8642 and n8895_not n8896_not ; n8898
g8643 and n8897_not n8898_not ; n8899
g8644 and b[44] n511 ; n8900
g8645 and b[42] n541 ; n8901
g8646 and b[43] n506 ; n8902
g8647 and n8901_not n8902_not ; n8903
g8648 and n8900_not n8903 ; n8904
g8649 and n514 n7072 ; n8905
g8650 and n8904 n8905_not ; n8906
g8651 and a[8] n8906_not ; n8907
g8652 and a[8] n8907_not ; n8908
g8653 and n8906_not n8907_not ; n8909
g8654 and n8908_not n8909_not ; n8910
g8655 and n8899 n8910_not ; n8911
g8656 and n8899_not n8910 ; n8912
g8657 and n8638_not n8912_not ; n8913
g8658 and n8911_not n8913 ; n8914
g8659 and n8638_not n8914_not ; n8915
g8660 and n8911_not n8914_not ; n8916
g8661 and n8912_not n8916 ; n8917
g8662 and n8915_not n8917_not ; n8918
g8663 and b[47] n362 ; n8919
g8664 and b[45] n403 ; n8920
g8665 and b[46] n357 ; n8921
g8666 and n8920_not n8921_not ; n8922
g8667 and n8919_not n8922 ; n8923
g8668 and n365 n7703 ; n8924
g8669 and n8923 n8924_not ; n8925
g8670 and a[5] n8925_not ; n8926
g8671 and a[5] n8926_not ; n8927
g8672 and n8925_not n8926_not ; n8928
g8673 and n8927_not n8928_not ; n8929
g8674 and n8918_not n8929_not ; n8930
g8675 and n8918_not n8930_not ; n8931
g8676 and n8929_not n8930_not ; n8932
g8677 and n8931_not n8932_not ; n8933
g8678 and n8606_not n8612_not ; n8934
g8679 and n8933 n8934 ; n8935
g8680 and n8933_not n8934_not ; n8936
g8681 and n8935_not n8936_not ; n8937
g8682 and b[50] n266 ; n8938
g8683 and b[48] n284 ; n8939
g8684 and b[49] n261 ; n8940
g8685 and n8939_not n8940_not ; n8941
g8686 and n8938_not n8941 ; n8942
g8687 and n8621_not n8623_not ; n8943
g8688 and b[49]_not b[50]_not ; n8944
g8689 and b[49] b[50] ; n8945
g8690 and n8944_not n8945_not ; n8946
g8691 and n8943_not n8946 ; n8947
g8692 and n8943 n8946_not ; n8948
g8693 and n8947_not n8948_not ; n8949
g8694 and n269 n8949 ; n8950
g8695 and n8942 n8950_not ; n8951
g8696 and a[2] n8951_not ; n8952
g8697 and a[2] n8952_not ; n8953
g8698 and n8951_not n8952_not ; n8954
g8699 and n8953_not n8954_not ; n8955
g8700 and n8937 n8955_not ; n8956
g8701 and n8937 n8956_not ; n8957
g8702 and n8955_not n8956_not ; n8958
g8703 and n8957_not n8958_not ; n8959
g8704 and n8633_not n8635_not ; n8960
g8705 and n8959_not n8960_not ; n8961
g8706 and n8959 n8960 ; n8962
g8707 and n8961_not n8962_not ; f[50]
g8708 and n8956_not n8961_not ; n8964
g8709 and b[51] n266 ; n8965
g8710 and b[49] n284 ; n8966
g8711 and b[50] n261 ; n8967
g8712 and n8966_not n8967_not ; n8968
g8713 and n8965_not n8968 ; n8969
g8714 and n8945_not n8947_not ; n8970
g8715 and b[50]_not b[51]_not ; n8971
g8716 and b[50] b[51] ; n8972
g8717 and n8971_not n8972_not ; n8973
g8718 and n8970_not n8973 ; n8974
g8719 and n8970 n8973_not ; n8975
g8720 and n8974_not n8975_not ; n8976
g8721 and n269 n8976 ; n8977
g8722 and n8969 n8977_not ; n8978
g8723 and a[2] n8978_not ; n8979
g8724 and a[2] n8979_not ; n8980
g8725 and n8978_not n8979_not ; n8981
g8726 and n8980_not n8981_not ; n8982
g8727 and n8930_not n8936_not ; n8983
g8728 and b[45] n511 ; n8984
g8729 and b[43] n541 ; n8985
g8730 and b[44] n506 ; n8986
g8731 and n8985_not n8986_not ; n8987
g8732 and n8984_not n8987 ; n8988
g8733 and n514 n7361 ; n8989
g8734 and n8988 n8989_not ; n8990
g8735 and a[8] n8990_not ; n8991
g8736 and a[8] n8991_not ; n8992
g8737 and n8990_not n8991_not ; n8993
g8738 and n8992_not n8993_not ; n8994
g8739 and n8854_not n8860_not ; n8995
g8740 and n8849_not n8851_not ; n8996
g8741 and b[33] n1627 ; n8997
g8742 and b[31] n1763 ; n8998
g8743 and b[32] n1622 ; n8999
g8744 and n8998_not n8999_not ; n9000
g8745 and n8997_not n9000 ; n9001
g8746 and n1630 n4223 ; n9002
g8747 and n9001 n9002_not ; n9003
g8748 and a[20] n9003_not ; n9004
g8749 and a[20] n9004_not ; n9005
g8750 and n9003_not n9004_not ; n9006
g8751 and n9005_not n9006_not ; n9007
g8752 and n8843_not n8845_not ; n9008
g8753 and n8837_not n8839_not ; n9009
g8754 and b[27] n2539 ; n9010
g8755 and b[25] n2685 ; n9011
g8756 and b[26] n2534 ; n9012
g8757 and n9011_not n9012_not ; n9013
g8758 and n9010_not n9013 ; n9014
g8759 and n2542 n2990 ; n9015
g8760 and n9014 n9015_not ; n9016
g8761 and a[26] n9016_not ; n9017
g8762 and a[26] n9017_not ; n9018
g8763 and n9016_not n9017_not ; n9019
g8764 and n9018_not n9019_not ; n9020
g8765 and n8779_not n8783_not ; n9021
g8766 and b[18] n4287 ; n9022
g8767 and b[16] n4532 ; n9023
g8768 and b[17] n4282 ; n9024
g8769 and n9023_not n9024_not ; n9025
g8770 and n9022_not n9025 ; n9026
g8771 and n1566 n4290 ; n9027
g8772 and n9026 n9027_not ; n9028
g8773 and a[35] n9028_not ; n9029
g8774 and a[35] n9029_not ; n9030
g8775 and n9028_not n9029_not ; n9031
g8776 and n9030_not n9031_not ; n9032
g8777 and n8772_not n8776_not ; n9033
g8778 and b[15] n5035 ; n9034
g8779 and b[13] n5277 ; n9035
g8780 and b[14] n5030 ; n9036
g8781 and n9035_not n9036_not ; n9037
g8782 and n9034_not n9037 ; n9038
g8783 and n1131 n5038 ; n9039
g8784 and n9038 n9039_not ; n9040
g8785 and a[38] n9040_not ; n9041
g8786 and a[38] n9041_not ; n9042
g8787 and n9040_not n9041_not ; n9043
g8788 and n9042_not n9043_not ; n9044
g8789 and n8767_not n8769_not ; n9045
g8790 and b[12] n5777 ; n9046
g8791 and b[10] n6059 ; n9047
g8792 and b[11] n5772 ; n9048
g8793 and n9047_not n9048_not ; n9049
g8794 and n9046_not n9049 ; n9050
g8795 and n842 n5780 ; n9051
g8796 and n9050 n9051_not ; n9052
g8797 and a[41] n9052_not ; n9053
g8798 and a[41] n9053_not ; n9054
g8799 and n9052_not n9053_not ; n9055
g8800 and n9054_not n9055_not ; n9056
g8801 and n8747_not n8751_not ; n9057
g8802 and b[6] n7446 ; n9058
g8803 and b[4] n7787 ; n9059
g8804 and b[5] n7441 ; n9060
g8805 and n9059_not n9060_not ; n9061
g8806 and n9058_not n9061 ; n9062
g8807 and n459 n7449 ; n9063
g8808 and n9062 n9063_not ; n9064
g8809 and a[47] n9064_not ; n9065
g8810 and a[47] n9065_not ; n9066
g8811 and n9064_not n9065_not ; n9067
g8812 and n9066_not n9067_not ; n9068
g8813 and a[50] a[51]_not ; n9069
g8814 and a[50]_not a[51] ; n9070
g8815 and n9069_not n9070_not ; n9071
g8816 and b[0] n9071_not ; n9072
g8817 and n8727_not n9072 ; n9073
g8818 and n8727 n9072_not ; n9074
g8819 and n9073_not n9074_not ; n9075
g8820 and b[3] n8362 ; n9076
g8821 and b[1] n8715 ; n9077
g8822 and b[2] n8357 ; n9078
g8823 and n9077_not n9078_not ; n9079
g8824 and n9076_not n9079 ; n9080
g8825 and n318 n8365 ; n9081
g8826 and n9080 n9081_not ; n9082
g8827 and a[50] n9082_not ; n9083
g8828 and a[50] n9083_not ; n9084
g8829 and n9082_not n9083_not ; n9085
g8830 and n9084_not n9085_not ; n9086
g8831 and n9075_not n9086_not ; n9087
g8832 and n9075 n9086 ; n9088
g8833 and n9087_not n9088_not ; n9089
g8834 and n9068_not n9089 ; n9090
g8835 and n9089 n9090_not ; n9091
g8836 and n9068_not n9090_not ; n9092
g8837 and n9091_not n9092_not ; n9093
g8838 and n8740_not n8744_not ; n9094
g8839 and n9093 n9094 ; n9095
g8840 and n9093_not n9094_not ; n9096
g8841 and n9095_not n9096_not ; n9097
g8842 and b[9] n6595 ; n9098
g8843 and b[7] n6902 ; n9099
g8844 and b[8] n6590 ; n9100
g8845 and n9099_not n9100_not ; n9101
g8846 and n9098_not n9101 ; n9102
g8847 and n651 n6598 ; n9103
g8848 and n9102 n9103_not ; n9104
g8849 and a[44] n9104_not ; n9105
g8850 and a[44] n9105_not ; n9106
g8851 and n9104_not n9105_not ; n9107
g8852 and n9106_not n9107_not ; n9108
g8853 and n9097_not n9108 ; n9109
g8854 and n9097 n9108_not ; n9110
g8855 and n9109_not n9110_not ; n9111
g8856 and n9057_not n9111 ; n9112
g8857 and n9057 n9111_not ; n9113
g8858 and n9112_not n9113_not ; n9114
g8859 and n9056_not n9114 ; n9115
g8860 and n9056_not n9115_not ; n9116
g8861 and n9114 n9115_not ; n9117
g8862 and n9116_not n9117_not ; n9118
g8863 and n9045_not n9118_not ; n9119
g8864 and n9045 n9117_not ; n9120
g8865 and n9116_not n9120 ; n9121
g8866 and n9119_not n9121_not ; n9122
g8867 and n9044_not n9122 ; n9123
g8868 and n9044 n9122_not ; n9124
g8869 and n9123_not n9124_not ; n9125
g8870 and n9033_not n9125 ; n9126
g8871 and n9033 n9125_not ; n9127
g8872 and n9126_not n9127_not ; n9128
g8873 and n9032_not n9128 ; n9129
g8874 and n9032 n9128_not ; n9130
g8875 and n9129_not n9130_not ; n9131
g8876 and n9021_not n9131 ; n9132
g8877 and n9021 n9131_not ; n9133
g8878 and n9132_not n9133_not ; n9134
g8879 and b[21] n3638 ; n9135
g8880 and b[19] n3843 ; n9136
g8881 and b[20] n3633 ; n9137
g8882 and n9136_not n9137_not ; n9138
g8883 and n9135_not n9138 ; n9139
g8884 and n1984 n3641 ; n9140
g8885 and n9139 n9140_not ; n9141
g8886 and a[32] n9141_not ; n9142
g8887 and a[32] n9142_not ; n9143
g8888 and n9141_not n9142_not ; n9144
g8889 and n9143_not n9144_not ; n9145
g8890 and n9134 n9145_not ; n9146
g8891 and n9134 n9146_not ; n9147
g8892 and n9145_not n9146_not ; n9148
g8893 and n9147_not n9148_not ; n9149
g8894 and n8798_not n8804_not ; n9150
g8895 and n9149 n9150 ; n9151
g8896 and n9149_not n9150_not ; n9152
g8897 and n9151_not n9152_not ; n9153
g8898 and b[24] n3050 ; n9154
g8899 and b[22] n3243 ; n9155
g8900 and b[23] n3045 ; n9156
g8901 and n9155_not n9156_not ; n9157
g8902 and n9154_not n9157 ; n9158
g8903 and n2458 n3053 ; n9159
g8904 and n9158 n9159_not ; n9160
g8905 and a[29] n9160_not ; n9161
g8906 and a[29] n9161_not ; n9162
g8907 and n9160_not n9161_not ; n9163
g8908 and n9162_not n9163_not ; n9164
g8909 and n9153_not n9164 ; n9165
g8910 and n9153 n9164_not ; n9166
g8911 and n9165_not n9166_not ; n9167
g8912 and n8822_not n9167 ; n9168
g8913 and n8822 n9167_not ; n9169
g8914 and n9168_not n9169_not ; n9170
g8915 and n9020_not n9170 ; n9171
g8916 and n9170 n9171_not ; n9172
g8917 and n9020_not n9171_not ; n9173
g8918 and n9172_not n9173_not ; n9174
g8919 and n9009_not n9174 ; n9175
g8920 and n9009 n9174_not ; n9176
g8921 and n9175_not n9176_not ; n9177
g8922 and b[30] n2048 ; n9178
g8923 and b[28] n2198 ; n9179
g8924 and b[29] n2043 ; n9180
g8925 and n9179_not n9180_not ; n9181
g8926 and n9178_not n9181 ; n9182
g8927 and n2051 n3577 ; n9183
g8928 and n9182 n9183_not ; n9184
g8929 and a[23] n9184_not ; n9185
g8930 and a[23] n9185_not ; n9186
g8931 and n9184_not n9185_not ; n9187
g8932 and n9186_not n9187_not ; n9188
g8933 and n9177_not n9188_not ; n9189
g8934 and n9177 n9188 ; n9190
g8935 and n9189_not n9190_not ; n9191
g8936 and n9008_not n9191 ; n9192
g8937 and n9008 n9191_not ; n9193
g8938 and n9192_not n9193_not ; n9194
g8939 and n9007_not n9194 ; n9195
g8940 and n9194 n9195_not ; n9196
g8941 and n9007_not n9195_not ; n9197
g8942 and n9196_not n9197_not ; n9198
g8943 and n8996_not n9198 ; n9199
g8944 and n8996 n9198_not ; n9200
g8945 and n9199_not n9200_not ; n9201
g8946 and b[36] n1302 ; n9202
g8947 and b[34] n1391 ; n9203
g8948 and b[35] n1297 ; n9204
g8949 and n9203_not n9204_not ; n9205
g8950 and n9202_not n9205 ; n9206
g8951 and n1305 n4922 ; n9207
g8952 and n9206 n9207_not ; n9208
g8953 and a[17] n9208_not ; n9209
g8954 and a[17] n9209_not ; n9210
g8955 and n9208_not n9209_not ; n9211
g8956 and n9210_not n9211_not ; n9212
g8957 and n9201_not n9212_not ; n9213
g8958 and n9201 n9212 ; n9214
g8959 and n9213_not n9214_not ; n9215
g8960 and n8995 n9215_not ; n9216
g8961 and n8995_not n9215 ; n9217
g8962 and n9216_not n9217_not ; n9218
g8963 and b[39] n951 ; n9219
g8964 and b[37] n1056 ; n9220
g8965 and b[38] n946 ; n9221
g8966 and n9220_not n9221_not ; n9222
g8967 and n9219_not n9222 ; n9223
g8968 and n954 n5451 ; n9224
g8969 and n9223 n9224_not ; n9225
g8970 and a[14] n9225_not ; n9226
g8971 and a[14] n9226_not ; n9227
g8972 and n9225_not n9226_not ; n9228
g8973 and n9227_not n9228_not ; n9229
g8974 and n9218 n9229_not ; n9230
g8975 and n9218 n9230_not ; n9231
g8976 and n9229_not n9230_not ; n9232
g8977 and n9231_not n9232_not ; n9233
g8978 and n8873_not n8879_not ; n9234
g8979 and n9233 n9234 ; n9235
g8980 and n9233_not n9234_not ; n9236
g8981 and n9235_not n9236_not ; n9237
g8982 and b[42] n700 ; n9238
g8983 and b[40] n767 ; n9239
g8984 and b[41] n695 ; n9240
g8985 and n9239_not n9240_not ; n9241
g8986 and n9238_not n9241 ; n9242
g8987 and n703 n6489 ; n9243
g8988 and n9242 n9243_not ; n9244
g8989 and a[11] n9244_not ; n9245
g8990 and a[11] n9245_not ; n9246
g8991 and n9244_not n9245_not ; n9247
g8992 and n9246_not n9247_not ; n9248
g8993 and n9237_not n9248 ; n9249
g8994 and n9237 n9248_not ; n9250
g8995 and n9249_not n9250_not ; n9251
g8996 and n8892_not n8898_not ; n9252
g8997 and n9251 n9252_not ; n9253
g8998 and n9251_not n9252 ; n9254
g8999 and n9253_not n9254_not ; n9255
g9000 and n8994_not n9255 ; n9256
g9001 and n9255 n9256_not ; n9257
g9002 and n8994_not n9256_not ; n9258
g9003 and n9257_not n9258_not ; n9259
g9004 and n8916_not n9259 ; n9260
g9005 and n8916 n9259_not ; n9261
g9006 and n9260_not n9261_not ; n9262
g9007 and b[48] n362 ; n9263
g9008 and b[46] n403 ; n9264
g9009 and b[47] n357 ; n9265
g9010 and n9264_not n9265_not ; n9266
g9011 and n9263_not n9266 ; n9267
g9012 and n365 n8009 ; n9268
g9013 and n9267 n9268_not ; n9269
g9014 and a[5] n9269_not ; n9270
g9015 and a[5] n9270_not ; n9271
g9016 and n9269_not n9270_not ; n9272
g9017 and n9271_not n9272_not ; n9273
g9018 and n9262 n9273 ; n9274
g9019 and n9262_not n9273_not ; n9275
g9020 and n9274_not n9275_not ; n9276
g9021 and n8983_not n9276 ; n9277
g9022 and n8983 n9276_not ; n9278
g9023 and n9277_not n9278_not ; n9279
g9024 and n8982_not n9279 ; n9280
g9025 and n8982 n9279_not ; n9281
g9026 and n9280_not n9281_not ; n9282
g9027 and n8964_not n9282 ; n9283
g9028 and n8964 n9282_not ; n9284
g9029 and n9283_not n9284_not ; f[51]
g9030 and n9280_not n9283_not ; n9286
g9031 and n9275_not n9277_not ; n9287
g9032 and n9250_not n9253_not ; n9288
g9033 and n9009_not n9174_not ; n9289
g9034 and n9171_not n9289_not ; n9290
g9035 and n9166_not n9168_not ; n9291
g9036 and n9129_not n9132_not ; n9292
g9037 and b[16] n5035 ; n9293
g9038 and b[14] n5277 ; n9294
g9039 and b[15] n5030 ; n9295
g9040 and n9294_not n9295_not ; n9296
g9041 and n9293_not n9296 ; n9297
g9042 and n1237 n5038 ; n9298
g9043 and n9297 n9298_not ; n9299
g9044 and a[38] n9299_not ; n9300
g9045 and a[38] n9300_not ; n9301
g9046 and n9299_not n9300_not ; n9302
g9047 and n9301_not n9302_not ; n9303
g9048 and n9115_not n9119_not ; n9304
g9049 and n9110_not n9112_not ; n9305
g9050 and b[7] n7446 ; n9306
g9051 and b[5] n7787 ; n9307
g9052 and b[6] n7441 ; n9308
g9053 and n9307_not n9308_not ; n9309
g9054 and n9306_not n9309 ; n9310
g9055 and n484 n7449 ; n9311
g9056 and n9310 n9311_not ; n9312
g9057 and a[47] n9312_not ; n9313
g9058 and a[47] n9313_not ; n9314
g9059 and n9312_not n9313_not ; n9315
g9060 and n9314_not n9315_not ; n9316
g9061 and n8727 n9072 ; n9317
g9062 and n9087_not n9317_not ; n9318
g9063 and b[4] n8362 ; n9319
g9064 and b[2] n8715 ; n9320
g9065 and b[3] n8357 ; n9321
g9066 and n9320_not n9321_not ; n9322
g9067 and n9319_not n9322 ; n9323
g9068 and n346 n8365 ; n9324
g9069 and n9323 n9324_not ; n9325
g9070 and a[50] n9325_not ; n9326
g9071 and a[50] n9326_not ; n9327
g9072 and n9325_not n9326_not ; n9328
g9073 and n9327_not n9328_not ; n9329
g9074 and a[53] n9072_not ; n9330
g9075 and a[51]_not a[52] ; n9331
g9076 and a[51] a[52]_not ; n9332
g9077 and n9331_not n9332_not ; n9333
g9078 and n9071 n9333_not ; n9334
g9079 and b[0] n9334 ; n9335
g9080 and a[52]_not a[53] ; n9336
g9081 and a[52] a[53]_not ; n9337
g9082 and n9336_not n9337_not ; n9338
g9083 and n9071_not n9338 ; n9339
g9084 and b[1] n9339 ; n9340
g9085 and n9335_not n9340_not ; n9341
g9086 and n9071_not n9338_not ; n9342
g9087 and n272_not n9342 ; n9343
g9088 and n9341 n9343_not ; n9344
g9089 and a[53] n9344_not ; n9345
g9090 and a[53] n9345_not ; n9346
g9091 and n9344_not n9345_not ; n9347
g9092 and n9346_not n9347_not ; n9348
g9093 and n9330 n9348_not ; n9349
g9094 and n9330_not n9348 ; n9350
g9095 and n9349_not n9350_not ; n9351
g9096 and n9329 n9351_not ; n9352
g9097 and n9329_not n9351 ; n9353
g9098 and n9352_not n9353_not ; n9354
g9099 and n9318_not n9354 ; n9355
g9100 and n9318 n9354_not ; n9356
g9101 and n9355_not n9356_not ; n9357
g9102 and n9316_not n9357 ; n9358
g9103 and n9357 n9358_not ; n9359
g9104 and n9316_not n9358_not ; n9360
g9105 and n9359_not n9360_not ; n9361
g9106 and n9090_not n9096_not ; n9362
g9107 and n9361 n9362 ; n9363
g9108 and n9361_not n9362_not ; n9364
g9109 and n9363_not n9364_not ; n9365
g9110 and b[10] n6595 ; n9366
g9111 and b[8] n6902 ; n9367
g9112 and b[9] n6590 ; n9368
g9113 and n9367_not n9368_not ; n9369
g9114 and n9366_not n9369 ; n9370
g9115 and n738 n6598 ; n9371
g9116 and n9370 n9371_not ; n9372
g9117 and a[44] n9372_not ; n9373
g9118 and a[44] n9373_not ; n9374
g9119 and n9372_not n9373_not ; n9375
g9120 and n9374_not n9375_not ; n9376
g9121 and n9365 n9376_not ; n9377
g9122 and n9365_not n9376 ; n9378
g9123 and n9305_not n9378_not ; n9379
g9124 and n9377_not n9379 ; n9380
g9125 and n9305_not n9380_not ; n9381
g9126 and n9377_not n9380_not ; n9382
g9127 and n9378_not n9382 ; n9383
g9128 and n9381_not n9383_not ; n9384
g9129 and b[13] n5777 ; n9385
g9130 and b[11] n6059 ; n9386
g9131 and b[12] n5772 ; n9387
g9132 and n9386_not n9387_not ; n9388
g9133 and n9385_not n9388 ; n9389
g9134 and n1008 n5780 ; n9390
g9135 and n9389 n9390_not ; n9391
g9136 and a[41] n9391_not ; n9392
g9137 and a[41] n9392_not ; n9393
g9138 and n9391_not n9392_not ; n9394
g9139 and n9393_not n9394_not ; n9395
g9140 and n9384 n9395 ; n9396
g9141 and n9384_not n9395_not ; n9397
g9142 and n9396_not n9397_not ; n9398
g9143 and n9304_not n9398 ; n9399
g9144 and n9304 n9398_not ; n9400
g9145 and n9399_not n9400_not ; n9401
g9146 and n9303_not n9401 ; n9402
g9147 and n9401 n9402_not ; n9403
g9148 and n9303_not n9402_not ; n9404
g9149 and n9403_not n9404_not ; n9405
g9150 and n9123_not n9126_not ; n9406
g9151 and n9405 n9406 ; n9407
g9152 and n9405_not n9406_not ; n9408
g9153 and n9407_not n9408_not ; n9409
g9154 and b[19] n4287 ; n9410
g9155 and b[17] n4532 ; n9411
g9156 and b[18] n4282 ; n9412
g9157 and n9411_not n9412_not ; n9413
g9158 and n9410_not n9413 ; n9414
g9159 and n1708 n4290 ; n9415
g9160 and n9414 n9415_not ; n9416
g9161 and a[35] n9416_not ; n9417
g9162 and a[35] n9417_not ; n9418
g9163 and n9416_not n9417_not ; n9419
g9164 and n9418_not n9419_not ; n9420
g9165 and n9409 n9420_not ; n9421
g9166 and n9409_not n9420 ; n9422
g9167 and n9292_not n9422_not ; n9423
g9168 and n9421_not n9423 ; n9424
g9169 and n9292_not n9424_not ; n9425
g9170 and n9421_not n9424_not ; n9426
g9171 and n9422_not n9426 ; n9427
g9172 and n9425_not n9427_not ; n9428
g9173 and b[22] n3638 ; n9429
g9174 and b[20] n3843 ; n9430
g9175 and b[21] n3633 ; n9431
g9176 and n9430_not n9431_not ; n9432
g9177 and n9429_not n9432 ; n9433
g9178 and n2145 n3641 ; n9434
g9179 and n9433 n9434_not ; n9435
g9180 and a[32] n9435_not ; n9436
g9181 and a[32] n9436_not ; n9437
g9182 and n9435_not n9436_not ; n9438
g9183 and n9437_not n9438_not ; n9439
g9184 and n9428_not n9439_not ; n9440
g9185 and n9428_not n9440_not ; n9441
g9186 and n9439_not n9440_not ; n9442
g9187 and n9441_not n9442_not ; n9443
g9188 and n9146_not n9152_not ; n9444
g9189 and n9443 n9444 ; n9445
g9190 and n9443_not n9444_not ; n9446
g9191 and n9445_not n9446_not ; n9447
g9192 and b[25] n3050 ; n9448
g9193 and b[23] n3243 ; n9449
g9194 and b[24] n3045 ; n9450
g9195 and n9449_not n9450_not ; n9451
g9196 and n9448_not n9451 ; n9452
g9197 and n2485 n3053 ; n9453
g9198 and n9452 n9453_not ; n9454
g9199 and a[29] n9454_not ; n9455
g9200 and a[29] n9455_not ; n9456
g9201 and n9454_not n9455_not ; n9457
g9202 and n9456_not n9457_not ; n9458
g9203 and n9447 n9458_not ; n9459
g9204 and n9447 n9459_not ; n9460
g9205 and n9458_not n9459_not ; n9461
g9206 and n9460_not n9461_not ; n9462
g9207 and n9291_not n9462 ; n9463
g9208 and n9291 n9462_not ; n9464
g9209 and n9463_not n9464_not ; n9465
g9210 and b[28] n2539 ; n9466
g9211 and b[26] n2685 ; n9467
g9212 and b[27] n2534 ; n9468
g9213 and n9467_not n9468_not ; n9469
g9214 and n9466_not n9469 ; n9470
g9215 and n2542 n3189 ; n9471
g9216 and n9470 n9471_not ; n9472
g9217 and a[26] n9472_not ; n9473
g9218 and a[26] n9473_not ; n9474
g9219 and n9472_not n9473_not ; n9475
g9220 and n9474_not n9475_not ; n9476
g9221 and n9465_not n9476_not ; n9477
g9222 and n9465 n9476 ; n9478
g9223 and n9477_not n9478_not ; n9479
g9224 and n9290 n9479_not ; n9480
g9225 and n9290_not n9479 ; n9481
g9226 and n9480_not n9481_not ; n9482
g9227 and b[31] n2048 ; n9483
g9228 and b[29] n2198 ; n9484
g9229 and b[30] n2043 ; n9485
g9230 and n9484_not n9485_not ; n9486
g9231 and n9483_not n9486 ; n9487
g9232 and n2051 n3796 ; n9488
g9233 and n9487 n9488_not ; n9489
g9234 and a[23] n9489_not ; n9490
g9235 and a[23] n9490_not ; n9491
g9236 and n9489_not n9490_not ; n9492
g9237 and n9491_not n9492_not ; n9493
g9238 and n9482 n9493_not ; n9494
g9239 and n9482 n9494_not ; n9495
g9240 and n9493_not n9494_not ; n9496
g9241 and n9495_not n9496_not ; n9497
g9242 and n9189_not n9192_not ; n9498
g9243 and n9497 n9498 ; n9499
g9244 and n9497_not n9498_not ; n9500
g9245 and n9499_not n9500_not ; n9501
g9246 and b[34] n1627 ; n9502
g9247 and b[32] n1763 ; n9503
g9248 and b[33] n1622 ; n9504
g9249 and n9503_not n9504_not ; n9505
g9250 and n9502_not n9505 ; n9506
g9251 and n1630 n4466 ; n9507
g9252 and n9506 n9507_not ; n9508
g9253 and a[20] n9508_not ; n9509
g9254 and a[20] n9509_not ; n9510
g9255 and n9508_not n9509_not ; n9511
g9256 and n9510_not n9511_not ; n9512
g9257 and n9501 n9512_not ; n9513
g9258 and n9501 n9513_not ; n9514
g9259 and n9512_not n9513_not ; n9515
g9260 and n9514_not n9515_not ; n9516
g9261 and n8996_not n9198_not ; n9517
g9262 and n9195_not n9517_not ; n9518
g9263 and n9516 n9518 ; n9519
g9264 and n9516_not n9518_not ; n9520
g9265 and n9519_not n9520_not ; n9521
g9266 and b[37] n1302 ; n9522
g9267 and b[35] n1391 ; n9523
g9268 and b[36] n1297 ; n9524
g9269 and n9523_not n9524_not ; n9525
g9270 and n9522_not n9525 ; n9526
g9271 and n1305 n5181 ; n9527
g9272 and n9526 n9527_not ; n9528
g9273 and a[17] n9528_not ; n9529
g9274 and a[17] n9529_not ; n9530
g9275 and n9528_not n9529_not ; n9531
g9276 and n9530_not n9531_not ; n9532
g9277 and n9521 n9532_not ; n9533
g9278 and n9521 n9533_not ; n9534
g9279 and n9532_not n9533_not ; n9535
g9280 and n9534_not n9535_not ; n9536
g9281 and n9213_not n9217_not ; n9537
g9282 and n9536 n9537 ; n9538
g9283 and n9536_not n9537_not ; n9539
g9284 and n9538_not n9539_not ; n9540
g9285 and b[40] n951 ; n9541
g9286 and b[38] n1056 ; n9542
g9287 and b[39] n946 ; n9543
g9288 and n9542_not n9543_not ; n9544
g9289 and n9541_not n9544 ; n9545
g9290 and n954 n5955 ; n9546
g9291 and n9545 n9546_not ; n9547
g9292 and a[14] n9547_not ; n9548
g9293 and a[14] n9548_not ; n9549
g9294 and n9547_not n9548_not ; n9550
g9295 and n9549_not n9550_not ; n9551
g9296 and n9540 n9551_not ; n9552
g9297 and n9540 n9552_not ; n9553
g9298 and n9551_not n9552_not ; n9554
g9299 and n9553_not n9554_not ; n9555
g9300 and n9230_not n9236_not ; n9556
g9301 and n9555 n9556 ; n9557
g9302 and n9555_not n9556_not ; n9558
g9303 and n9557_not n9558_not ; n9559
g9304 and b[43] n700 ; n9560
g9305 and b[41] n767 ; n9561
g9306 and b[42] n695 ; n9562
g9307 and n9561_not n9562_not ; n9563
g9308 and n9560_not n9563 ; n9564
g9309 and n703 n6515 ; n9565
g9310 and n9564 n9565_not ; n9566
g9311 and a[11] n9566_not ; n9567
g9312 and a[11] n9567_not ; n9568
g9313 and n9566_not n9567_not ; n9569
g9314 and n9568_not n9569_not ; n9570
g9315 and n9559 n9570_not ; n9571
g9316 and n9559_not n9570 ; n9572
g9317 and n9288_not n9572_not ; n9573
g9318 and n9571_not n9573 ; n9574
g9319 and n9288_not n9574_not ; n9575
g9320 and n9571_not n9574_not ; n9576
g9321 and n9572_not n9576 ; n9577
g9322 and n9575_not n9577_not ; n9578
g9323 and b[46] n511 ; n9579
g9324 and b[44] n541 ; n9580
g9325 and b[45] n506 ; n9581
g9326 and n9580_not n9581_not ; n9582
g9327 and n9579_not n9582 ; n9583
g9328 and n514 n7677 ; n9584
g9329 and n9583 n9584_not ; n9585
g9330 and a[8] n9585_not ; n9586
g9331 and a[8] n9586_not ; n9587
g9332 and n9585_not n9586_not ; n9588
g9333 and n9587_not n9588_not ; n9589
g9334 and n9578_not n9589_not ; n9590
g9335 and n9578_not n9590_not ; n9591
g9336 and n9589_not n9590_not ; n9592
g9337 and n9591_not n9592_not ; n9593
g9338 and n8916_not n9259_not ; n9594
g9339 and n9256_not n9594_not ; n9595
g9340 and n9593 n9595 ; n9596
g9341 and n9593_not n9595_not ; n9597
g9342 and n9596_not n9597_not ; n9598
g9343 and b[49] n362 ; n9599
g9344 and b[47] n403 ; n9600
g9345 and b[48] n357 ; n9601
g9346 and n9600_not n9601_not ; n9602
g9347 and n9599_not n9602 ; n9603
g9348 and n365 n8625 ; n9604
g9349 and n9603 n9604_not ; n9605
g9350 and a[5] n9605_not ; n9606
g9351 and a[5] n9606_not ; n9607
g9352 and n9605_not n9606_not ; n9608
g9353 and n9607_not n9608_not ; n9609
g9354 and n9598 n9609_not ; n9610
g9355 and n9598 n9610_not ; n9611
g9356 and n9609_not n9610_not ; n9612
g9357 and n9611_not n9612_not ; n9613
g9358 and n9287_not n9613 ; n9614
g9359 and n9287 n9613_not ; n9615
g9360 and n9614_not n9615_not ; n9616
g9361 and b[52] n266 ; n9617
g9362 and b[50] n284 ; n9618
g9363 and b[51] n261 ; n9619
g9364 and n9618_not n9619_not ; n9620
g9365 and n9617_not n9620 ; n9621
g9366 and n8972_not n8974_not ; n9622
g9367 and b[51]_not b[52]_not ; n9623
g9368 and b[51] b[52] ; n9624
g9369 and n9623_not n9624_not ; n9625
g9370 and n9622_not n9625 ; n9626
g9371 and n9622 n9625_not ; n9627
g9372 and n9626_not n9627_not ; n9628
g9373 and n269 n9628 ; n9629
g9374 and n9621 n9629_not ; n9630
g9375 and a[2] n9630_not ; n9631
g9376 and a[2] n9631_not ; n9632
g9377 and n9630_not n9631_not ; n9633
g9378 and n9632_not n9633_not ; n9634
g9379 and n9616_not n9634_not ; n9635
g9380 and n9616 n9634 ; n9636
g9381 and n9635_not n9636_not ; n9637
g9382 and n9286_not n9637 ; n9638
g9383 and n9286 n9637_not ; n9639
g9384 and n9638_not n9639_not ; f[52]
g9385 and n9635_not n9638_not ; n9641
g9386 and n9287_not n9613_not ; n9642
g9387 and n9610_not n9642_not ; n9643
g9388 and b[35] n1627 ; n9644
g9389 and b[33] n1763 ; n9645
g9390 and b[34] n1622 ; n9646
g9391 and n9645_not n9646_not ; n9647
g9392 and n9644_not n9647 ; n9648
g9393 and n1630 n4696 ; n9649
g9394 and n9648 n9649_not ; n9650
g9395 and a[20] n9650_not ; n9651
g9396 and a[20] n9651_not ; n9652
g9397 and n9650_not n9651_not ; n9653
g9398 and n9652_not n9653_not ; n9654
g9399 and n9494_not n9500_not ; n9655
g9400 and b[32] n2048 ; n9656
g9401 and b[30] n2198 ; n9657
g9402 and b[31] n2043 ; n9658
g9403 and n9657_not n9658_not ; n9659
g9404 and n9656_not n9659 ; n9660
g9405 and n2051 n4013 ; n9661
g9406 and n9660 n9661_not ; n9662
g9407 and a[23] n9662_not ; n9663
g9408 and a[23] n9663_not ; n9664
g9409 and n9662_not n9663_not ; n9665
g9410 and n9664_not n9665_not ; n9666
g9411 and n9477_not n9481_not ; n9667
g9412 and b[29] n2539 ; n9668
g9413 and b[27] n2685 ; n9669
g9414 and b[28] n2534 ; n9670
g9415 and n9669_not n9670_not ; n9671
g9416 and n9668_not n9671 ; n9672
g9417 and n2542 n3383 ; n9673
g9418 and n9672 n9673_not ; n9674
g9419 and a[26] n9674_not ; n9675
g9420 and a[26] n9675_not ; n9676
g9421 and n9674_not n9675_not ; n9677
g9422 and n9676_not n9677_not ; n9678
g9423 and n9291_not n9462_not ; n9679
g9424 and n9459_not n9679_not ; n9680
g9425 and n9440_not n9446_not ; n9681
g9426 and b[23] n3638 ; n9682
g9427 and b[21] n3843 ; n9683
g9428 and b[22] n3633 ; n9684
g9429 and n9683_not n9684_not ; n9685
g9430 and n9682_not n9685 ; n9686
g9431 and n2300 n3641 ; n9687
g9432 and n9686 n9687_not ; n9688
g9433 and a[32] n9688_not ; n9689
g9434 and a[32] n9689_not ; n9690
g9435 and n9688_not n9689_not ; n9691
g9436 and n9690_not n9691_not ; n9692
g9437 and n9402_not n9408_not ; n9693
g9438 and b[17] n5035 ; n9694
g9439 and b[15] n5277 ; n9695
g9440 and b[16] n5030 ; n9696
g9441 and n9695_not n9696_not ; n9697
g9442 and n9694_not n9697 ; n9698
g9443 and n1356 n5038 ; n9699
g9444 and n9698 n9699_not ; n9700
g9445 and a[38] n9700_not ; n9701
g9446 and a[38] n9701_not ; n9702
g9447 and n9700_not n9701_not ; n9703
g9448 and n9702_not n9703_not ; n9704
g9449 and n9397_not n9399_not ; n9705
g9450 and b[14] n5777 ; n9706
g9451 and b[12] n6059 ; n9707
g9452 and b[13] n5772 ; n9708
g9453 and n9707_not n9708_not ; n9709
g9454 and n9706_not n9709 ; n9710
g9455 and n1034 n5780 ; n9711
g9456 and n9710 n9711_not ; n9712
g9457 and a[41] n9712_not ; n9713
g9458 and a[41] n9713_not ; n9714
g9459 and n9712_not n9713_not ; n9715
g9460 and n9714_not n9715_not ; n9716
g9461 and b[11] n6595 ; n9717
g9462 and b[9] n6902 ; n9718
g9463 and b[10] n6590 ; n9719
g9464 and n9718_not n9719_not ; n9720
g9465 and n9717_not n9720 ; n9721
g9466 and n818 n6598 ; n9722
g9467 and n9721 n9722_not ; n9723
g9468 and a[44] n9723_not ; n9724
g9469 and a[44] n9724_not ; n9725
g9470 and n9723_not n9724_not ; n9726
g9471 and n9725_not n9726_not ; n9727
g9472 and n9358_not n9364_not ; n9728
g9473 and n9353_not n9355_not ; n9729
g9474 and b[2] n9339 ; n9730
g9475 and n9071 n9338_not ; n9731
g9476 and n9333 n9731 ; n9732
g9477 and b[0] n9732 ; n9733
g9478 and b[1] n9334 ; n9734
g9479 and n9733_not n9734_not ; n9735
g9480 and n9730_not n9735 ; n9736
g9481 and n296 n9342 ; n9737
g9482 and n9736 n9737_not ; n9738
g9483 and a[53] n9738_not ; n9739
g9484 and a[53] n9739_not ; n9740
g9485 and n9738_not n9739_not ; n9741
g9486 and n9740_not n9741_not ; n9742
g9487 and n9349_not n9742 ; n9743
g9488 and n9349 n9742_not ; n9744
g9489 and n9743_not n9744_not ; n9745
g9490 and b[5] n8362 ; n9746
g9491 and b[3] n8715 ; n9747
g9492 and b[4] n8357 ; n9748
g9493 and n9747_not n9748_not ; n9749
g9494 and n9746_not n9749 ; n9750
g9495 and n394 n8365 ; n9751
g9496 and n9750 n9751_not ; n9752
g9497 and a[50] n9752_not ; n9753
g9498 and a[50] n9753_not ; n9754
g9499 and n9752_not n9753_not ; n9755
g9500 and n9754_not n9755_not ; n9756
g9501 and n9745 n9756_not ; n9757
g9502 and n9745_not n9756 ; n9758
g9503 and n9729_not n9758_not ; n9759
g9504 and n9757_not n9759 ; n9760
g9505 and n9729_not n9760_not ; n9761
g9506 and n9757_not n9760_not ; n9762
g9507 and n9758_not n9762 ; n9763
g9508 and n9761_not n9763_not ; n9764
g9509 and b[8] n7446 ; n9765
g9510 and b[6] n7787 ; n9766
g9511 and b[7] n7441 ; n9767
g9512 and n9766_not n9767_not ; n9768
g9513 and n9765_not n9768 ; n9769
g9514 and n585 n7449 ; n9770
g9515 and n9769 n9770_not ; n9771
g9516 and a[47] n9771_not ; n9772
g9517 and a[47] n9772_not ; n9773
g9518 and n9771_not n9772_not ; n9774
g9519 and n9773_not n9774_not ; n9775
g9520 and n9764 n9775 ; n9776
g9521 and n9764_not n9775_not ; n9777
g9522 and n9776_not n9777_not ; n9778
g9523 and n9728_not n9778 ; n9779
g9524 and n9728 n9778_not ; n9780
g9525 and n9779_not n9780_not ; n9781
g9526 and n9727 n9781_not ; n9782
g9527 and n9727_not n9781 ; n9783
g9528 and n9782_not n9783_not ; n9784
g9529 and n9382_not n9784 ; n9785
g9530 and n9382 n9784_not ; n9786
g9531 and n9785_not n9786_not ; n9787
g9532 and n9716_not n9787 ; n9788
g9533 and n9787 n9788_not ; n9789
g9534 and n9716_not n9788_not ; n9790
g9535 and n9789_not n9790_not ; n9791
g9536 and n9705_not n9791_not ; n9792
g9537 and n9705 n9791 ; n9793
g9538 and n9792_not n9793_not ; n9794
g9539 and n9704_not n9794 ; n9795
g9540 and n9704_not n9795_not ; n9796
g9541 and n9794 n9795_not ; n9797
g9542 and n9796_not n9797_not ; n9798
g9543 and n9693_not n9798_not ; n9799
g9544 and n9693_not n9799_not ; n9800
g9545 and n9798_not n9799_not ; n9801
g9546 and n9800_not n9801_not ; n9802
g9547 and b[20] n4287 ; n9803
g9548 and b[18] n4532 ; n9804
g9549 and b[19] n4282 ; n9805
g9550 and n9804_not n9805_not ; n9806
g9551 and n9803_not n9806 ; n9807
g9552 and n1846 n4290 ; n9808
g9553 and n9807 n9808_not ; n9809
g9554 and a[35] n9809_not ; n9810
g9555 and a[35] n9810_not ; n9811
g9556 and n9809_not n9810_not ; n9812
g9557 and n9811_not n9812_not ; n9813
g9558 and n9802_not n9813_not ; n9814
g9559 and n9802_not n9814_not ; n9815
g9560 and n9813_not n9814_not ; n9816
g9561 and n9815_not n9816_not ; n9817
g9562 and n9426_not n9817_not ; n9818
g9563 and n9426 n9817 ; n9819
g9564 and n9818_not n9819_not ; n9820
g9565 and n9692_not n9820 ; n9821
g9566 and n9692_not n9821_not ; n9822
g9567 and n9820 n9821_not ; n9823
g9568 and n9822_not n9823_not ; n9824
g9569 and n9681_not n9824_not ; n9825
g9570 and n9681_not n9825_not ; n9826
g9571 and n9824_not n9825_not ; n9827
g9572 and n9826_not n9827_not ; n9828
g9573 and b[26] n3050 ; n9829
g9574 and b[24] n3243 ; n9830
g9575 and b[25] n3045 ; n9831
g9576 and n9830_not n9831_not ; n9832
g9577 and n9829_not n9832 ; n9833
g9578 and n2813 n3053 ; n9834
g9579 and n9833 n9834_not ; n9835
g9580 and a[29] n9835_not ; n9836
g9581 and a[29] n9836_not ; n9837
g9582 and n9835_not n9836_not ; n9838
g9583 and n9837_not n9838_not ; n9839
g9584 and n9828 n9839 ; n9840
g9585 and n9828_not n9839_not ; n9841
g9586 and n9840_not n9841_not ; n9842
g9587 and n9680_not n9842 ; n9843
g9588 and n9680 n9842_not ; n9844
g9589 and n9843_not n9844_not ; n9845
g9590 and n9678 n9845_not ; n9846
g9591 and n9678_not n9845 ; n9847
g9592 and n9846_not n9847_not ; n9848
g9593 and n9667_not n9848 ; n9849
g9594 and n9667 n9848_not ; n9850
g9595 and n9849_not n9850_not ; n9851
g9596 and n9666 n9851_not ; n9852
g9597 and n9666_not n9851 ; n9853
g9598 and n9852_not n9853_not ; n9854
g9599 and n9655_not n9854 ; n9855
g9600 and n9655 n9854_not ; n9856
g9601 and n9855_not n9856_not ; n9857
g9602 and n9654_not n9857 ; n9858
g9603 and n9857 n9858_not ; n9859
g9604 and n9654_not n9858_not ; n9860
g9605 and n9859_not n9860_not ; n9861
g9606 and n9513_not n9520_not ; n9862
g9607 and n9861 n9862 ; n9863
g9608 and n9861_not n9862_not ; n9864
g9609 and n9863_not n9864_not ; n9865
g9610 and b[38] n1302 ; n9866
g9611 and b[36] n1391 ; n9867
g9612 and b[37] n1297 ; n9868
g9613 and n9867_not n9868_not ; n9869
g9614 and n9866_not n9869 ; n9870
g9615 and n1305 n5205 ; n9871
g9616 and n9870 n9871_not ; n9872
g9617 and a[17] n9872_not ; n9873
g9618 and a[17] n9873_not ; n9874
g9619 and n9872_not n9873_not ; n9875
g9620 and n9874_not n9875_not ; n9876
g9621 and n9865 n9876_not ; n9877
g9622 and n9865 n9877_not ; n9878
g9623 and n9876_not n9877_not ; n9879
g9624 and n9878_not n9879_not ; n9880
g9625 and n9533_not n9539_not ; n9881
g9626 and n9880 n9881 ; n9882
g9627 and n9880_not n9881_not ; n9883
g9628 and n9882_not n9883_not ; n9884
g9629 and b[41] n951 ; n9885
g9630 and b[39] n1056 ; n9886
g9631 and b[40] n946 ; n9887
g9632 and n9886_not n9887_not ; n9888
g9633 and n9885_not n9888 ; n9889
g9634 and n954 n6219 ; n9890
g9635 and n9889 n9890_not ; n9891
g9636 and a[14] n9891_not ; n9892
g9637 and a[14] n9892_not ; n9893
g9638 and n9891_not n9892_not ; n9894
g9639 and n9893_not n9894_not ; n9895
g9640 and n9884 n9895_not ; n9896
g9641 and n9884 n9896_not ; n9897
g9642 and n9895_not n9896_not ; n9898
g9643 and n9897_not n9898_not ; n9899
g9644 and n9552_not n9558_not ; n9900
g9645 and n9899 n9900 ; n9901
g9646 and n9899_not n9900_not ; n9902
g9647 and n9901_not n9902_not ; n9903
g9648 and b[44] n700 ; n9904
g9649 and b[42] n767 ; n9905
g9650 and b[43] n695 ; n9906
g9651 and n9905_not n9906_not ; n9907
g9652 and n9904_not n9907 ; n9908
g9653 and n703 n7072 ; n9909
g9654 and n9908 n9909_not ; n9910
g9655 and a[11] n9910_not ; n9911
g9656 and a[11] n9911_not ; n9912
g9657 and n9910_not n9911_not ; n9913
g9658 and n9912_not n9913_not ; n9914
g9659 and n9903 n9914_not ; n9915
g9660 and n9903_not n9914 ; n9916
g9661 and n9576_not n9916_not ; n9917
g9662 and n9915_not n9917 ; n9918
g9663 and n9576_not n9918_not ; n9919
g9664 and n9915_not n9918_not ; n9920
g9665 and n9916_not n9920 ; n9921
g9666 and n9919_not n9921_not ; n9922
g9667 and b[47] n511 ; n9923
g9668 and b[45] n541 ; n9924
g9669 and b[46] n506 ; n9925
g9670 and n9924_not n9925_not ; n9926
g9671 and n9923_not n9926 ; n9927
g9672 and n514 n7703 ; n9928
g9673 and n9927 n9928_not ; n9929
g9674 and a[8] n9929_not ; n9930
g9675 and a[8] n9930_not ; n9931
g9676 and n9929_not n9930_not ; n9932
g9677 and n9931_not n9932_not ; n9933
g9678 and n9922_not n9933_not ; n9934
g9679 and n9922_not n9934_not ; n9935
g9680 and n9933_not n9934_not ; n9936
g9681 and n9935_not n9936_not ; n9937
g9682 and n9590_not n9597_not ; n9938
g9683 and n9937 n9938 ; n9939
g9684 and n9937_not n9938_not ; n9940
g9685 and n9939_not n9940_not ; n9941
g9686 and b[50] n362 ; n9942
g9687 and b[48] n403 ; n9943
g9688 and b[49] n357 ; n9944
g9689 and n9943_not n9944_not ; n9945
g9690 and n9942_not n9945 ; n9946
g9691 and n365 n8949 ; n9947
g9692 and n9946 n9947_not ; n9948
g9693 and a[5] n9948_not ; n9949
g9694 and a[5] n9949_not ; n9950
g9695 and n9948_not n9949_not ; n9951
g9696 and n9950_not n9951_not ; n9952
g9697 and n9941 n9952_not ; n9953
g9698 and n9941_not n9952 ; n9954
g9699 and n9643_not n9954_not ; n9955
g9700 and n9953_not n9955 ; n9956
g9701 and n9643_not n9956_not ; n9957
g9702 and n9953_not n9956_not ; n9958
g9703 and n9954_not n9958 ; n9959
g9704 and n9957_not n9959_not ; n9960
g9705 and b[53] n266 ; n9961
g9706 and b[51] n284 ; n9962
g9707 and b[52] n261 ; n9963
g9708 and n9962_not n9963_not ; n9964
g9709 and n9961_not n9964 ; n9965
g9710 and n9624_not n9626_not ; n9966
g9711 and b[52]_not b[53]_not ; n9967
g9712 and b[52] b[53] ; n9968
g9713 and n9967_not n9968_not ; n9969
g9714 and n9966_not n9969 ; n9970
g9715 and n9966 n9969_not ; n9971
g9716 and n9970_not n9971_not ; n9972
g9717 and n269 n9972 ; n9973
g9718 and n9965 n9973_not ; n9974
g9719 and a[2] n9974_not ; n9975
g9720 and a[2] n9975_not ; n9976
g9721 and n9974_not n9975_not ; n9977
g9722 and n9976_not n9977_not ; n9978
g9723 and n9960_not n9978 ; n9979
g9724 and n9960 n9978_not ; n9980
g9725 and n9979_not n9980_not ; n9981
g9726 and n9641_not n9981_not ; n9982
g9727 and n9641 n9981 ; n9983
g9728 and n9982_not n9983_not ; f[53]
g9729 and n9960_not n9978_not ; n9985
g9730 and n9982_not n9985_not ; n9986
g9731 and b[54] n266 ; n9987
g9732 and b[52] n284 ; n9988
g9733 and b[53] n261 ; n9989
g9734 and n9988_not n9989_not ; n9990
g9735 and n9987_not n9990 ; n9991
g9736 and n9968_not n9970_not ; n9992
g9737 and b[53]_not b[54]_not ; n9993
g9738 and b[53] b[54] ; n9994
g9739 and n9993_not n9994_not ; n9995
g9740 and n9992_not n9995 ; n9996
g9741 and n9992 n9995_not ; n9997
g9742 and n9996_not n9997_not ; n9998
g9743 and n269 n9998 ; n9999
g9744 and n9991 n9999_not ; n10000
g9745 and a[2] n10000_not ; n10001
g9746 and a[2] n10001_not ; n10002
g9747 and n10000_not n10001_not ; n10003
g9748 and n10002_not n10003_not ; n10004
g9749 and b[45] n700 ; n10005
g9750 and b[43] n767 ; n10006
g9751 and b[44] n695 ; n10007
g9752 and n10006_not n10007_not ; n10008
g9753 and n10005_not n10008 ; n10009
g9754 and n703 n7361 ; n10010
g9755 and n10009 n10010_not ; n10011
g9756 and a[11] n10011_not ; n10012
g9757 and a[11] n10012_not ; n10013
g9758 and n10011_not n10012_not ; n10014
g9759 and n10013_not n10014_not ; n10015
g9760 and n9896_not n9902_not ; n10016
g9761 and n9858_not n9864_not ; n10017
g9762 and n9853_not n9855_not ; n10018
g9763 and n9847_not n9849_not ; n10019
g9764 and b[30] n2539 ; n10020
g9765 and b[28] n2685 ; n10021
g9766 and b[29] n2534 ; n10022
g9767 and n10021_not n10022_not ; n10023
g9768 and n10020_not n10023 ; n10024
g9769 and n2542 n3577 ; n10025
g9770 and n10024 n10025_not ; n10026
g9771 and a[26] n10026_not ; n10027
g9772 and a[26] n10027_not ; n10028
g9773 and n10026_not n10027_not ; n10029
g9774 and n10028_not n10029_not ; n10030
g9775 and n9841_not n9843_not ; n10031
g9776 and b[27] n3050 ; n10032
g9777 and b[25] n3243 ; n10033
g9778 and b[26] n3045 ; n10034
g9779 and n10033_not n10034_not ; n10035
g9780 and n10032_not n10035 ; n10036
g9781 and n2990 n3053 ; n10037
g9782 and n10036 n10037_not ; n10038
g9783 and a[29] n10038_not ; n10039
g9784 and a[29] n10039_not ; n10040
g9785 and n10038_not n10039_not ; n10041
g9786 and n10040_not n10041_not ; n10042
g9787 and n9821_not n9825_not ; n10043
g9788 and b[24] n3638 ; n10044
g9789 and b[22] n3843 ; n10045
g9790 and b[23] n3633 ; n10046
g9791 and n10045_not n10046_not ; n10047
g9792 and n10044_not n10047 ; n10048
g9793 and n2458 n3641 ; n10049
g9794 and n10048 n10049_not ; n10050
g9795 and a[32] n10050_not ; n10051
g9796 and a[32] n10051_not ; n10052
g9797 and n10050_not n10051_not ; n10053
g9798 and n10052_not n10053_not ; n10054
g9799 and n9814_not n9818_not ; n10055
g9800 and b[21] n4287 ; n10056
g9801 and b[19] n4532 ; n10057
g9802 and b[20] n4282 ; n10058
g9803 and n10057_not n10058_not ; n10059
g9804 and n10056_not n10059 ; n10060
g9805 and n1984 n4290 ; n10061
g9806 and n10060 n10061_not ; n10062
g9807 and a[35] n10062_not ; n10063
g9808 and a[35] n10063_not ; n10064
g9809 and n10062_not n10063_not ; n10065
g9810 and n10064_not n10065_not ; n10066
g9811 and n9795_not n9799_not ; n10067
g9812 and b[18] n5035 ; n10068
g9813 and b[16] n5277 ; n10069
g9814 and b[17] n5030 ; n10070
g9815 and n10069_not n10070_not ; n10071
g9816 and n10068_not n10071 ; n10072
g9817 and n1566 n5038 ; n10073
g9818 and n10072 n10073_not ; n10074
g9819 and a[38] n10074_not ; n10075
g9820 and a[38] n10075_not ; n10076
g9821 and n10074_not n10075_not ; n10077
g9822 and n10076_not n10077_not ; n10078
g9823 and n9788_not n9792_not ; n10079
g9824 and b[15] n5777 ; n10080
g9825 and b[13] n6059 ; n10081
g9826 and b[14] n5772 ; n10082
g9827 and n10081_not n10082_not ; n10083
g9828 and n10080_not n10083 ; n10084
g9829 and n1131 n5780 ; n10085
g9830 and n10084 n10085_not ; n10086
g9831 and a[41] n10086_not ; n10087
g9832 and a[41] n10087_not ; n10088
g9833 and n10086_not n10087_not ; n10089
g9834 and n10088_not n10089_not ; n10090
g9835 and n9783_not n9785_not ; n10091
g9836 and b[12] n6595 ; n10092
g9837 and b[10] n6902 ; n10093
g9838 and b[11] n6590 ; n10094
g9839 and n10093_not n10094_not ; n10095
g9840 and n10092_not n10095 ; n10096
g9841 and n842 n6598 ; n10097
g9842 and n10096 n10097_not ; n10098
g9843 and a[44] n10098_not ; n10099
g9844 and a[44] n10099_not ; n10100
g9845 and n10098_not n10099_not ; n10101
g9846 and n10100_not n10101_not ; n10102
g9847 and n9777_not n9779_not ; n10103
g9848 and b[9] n7446 ; n10104
g9849 and b[7] n7787 ; n10105
g9850 and b[8] n7441 ; n10106
g9851 and n10105_not n10106_not ; n10107
g9852 and n10104_not n10107 ; n10108
g9853 and n651 n7449 ; n10109
g9854 and n10108 n10109_not ; n10110
g9855 and a[47] n10110_not ; n10111
g9856 and a[47] n10111_not ; n10112
g9857 and n10110_not n10111_not ; n10113
g9858 and n10112_not n10113_not ; n10114
g9859 and b[6] n8362 ; n10115
g9860 and b[4] n8715 ; n10116
g9861 and b[5] n8357 ; n10117
g9862 and n10116_not n10117_not ; n10118
g9863 and n10115_not n10118 ; n10119
g9864 and n459 n8365 ; n10120
g9865 and n10119 n10120_not ; n10121
g9866 and a[50] n10121_not ; n10122
g9867 and a[50] n10122_not ; n10123
g9868 and n10121_not n10122_not ; n10124
g9869 and n10123_not n10124_not ; n10125
g9870 and a[53] a[54]_not ; n10126
g9871 and a[53]_not a[54] ; n10127
g9872 and n10126_not n10127_not ; n10128
g9873 and b[0] n10128_not ; n10129
g9874 and n9744_not n10129 ; n10130
g9875 and n9744 n10129_not ; n10131
g9876 and n10130_not n10131_not ; n10132
g9877 and b[3] n9339 ; n10133
g9878 and b[1] n9732 ; n10134
g9879 and b[2] n9334 ; n10135
g9880 and n10134_not n10135_not ; n10136
g9881 and n10133_not n10136 ; n10137
g9882 and n318 n9342 ; n10138
g9883 and n10137 n10138_not ; n10139
g9884 and a[53] n10139_not ; n10140
g9885 and a[53] n10140_not ; n10141
g9886 and n10139_not n10140_not ; n10142
g9887 and n10141_not n10142_not ; n10143
g9888 and n10132_not n10143_not ; n10144
g9889 and n10132 n10143 ; n10145
g9890 and n10144_not n10145_not ; n10146
g9891 and n10125_not n10146 ; n10147
g9892 and n10146 n10147_not ; n10148
g9893 and n10125_not n10147_not ; n10149
g9894 and n10148_not n10149_not ; n10150
g9895 and n9762_not n10150_not ; n10151
g9896 and n9762 n10150 ; n10152
g9897 and n10151_not n10152_not ; n10153
g9898 and n10114_not n10153 ; n10154
g9899 and n10114_not n10154_not ; n10155
g9900 and n10153 n10154_not ; n10156
g9901 and n10155_not n10156_not ; n10157
g9902 and n10103_not n10157_not ; n10158
g9903 and n10103 n10156_not ; n10159
g9904 and n10155_not n10159 ; n10160
g9905 and n10158_not n10160_not ; n10161
g9906 and n10102_not n10161 ; n10162
g9907 and n10102_not n10162_not ; n10163
g9908 and n10161 n10162_not ; n10164
g9909 and n10163_not n10164_not ; n10165
g9910 and n10091_not n10165_not ; n10166
g9911 and n10091 n10164_not ; n10167
g9912 and n10163_not n10167 ; n10168
g9913 and n10166_not n10168_not ; n10169
g9914 and n10090_not n10169 ; n10170
g9915 and n10090 n10169_not ; n10171
g9916 and n10170_not n10171_not ; n10172
g9917 and n10079_not n10172 ; n10173
g9918 and n10079 n10172_not ; n10174
g9919 and n10173_not n10174_not ; n10175
g9920 and n10078_not n10175 ; n10176
g9921 and n10078_not n10176_not ; n10177
g9922 and n10175 n10176_not ; n10178
g9923 and n10177_not n10178_not ; n10179
g9924 and n10067_not n10179_not ; n10180
g9925 and n10067 n10178_not ; n10181
g9926 and n10177_not n10181 ; n10182
g9927 and n10180_not n10182_not ; n10183
g9928 and n10066_not n10183 ; n10184
g9929 and n10066 n10183_not ; n10185
g9930 and n10184_not n10185_not ; n10186
g9931 and n10055_not n10186 ; n10187
g9932 and n10055 n10186_not ; n10188
g9933 and n10187_not n10188_not ; n10189
g9934 and n10054_not n10189 ; n10190
g9935 and n10054 n10189_not ; n10191
g9936 and n10190_not n10191_not ; n10192
g9937 and n10043_not n10192 ; n10193
g9938 and n10043 n10192_not ; n10194
g9939 and n10193_not n10194_not ; n10195
g9940 and n10042_not n10195 ; n10196
g9941 and n10042 n10195_not ; n10197
g9942 and n10196_not n10197_not ; n10198
g9943 and n10031_not n10198 ; n10199
g9944 and n10031 n10198_not ; n10200
g9945 and n10199_not n10200_not ; n10201
g9946 and n10030_not n10201 ; n10202
g9947 and n10030 n10201_not ; n10203
g9948 and n10202_not n10203_not ; n10204
g9949 and n10019_not n10204 ; n10205
g9950 and n10019 n10204_not ; n10206
g9951 and n10205_not n10206_not ; n10207
g9952 and b[33] n2048 ; n10208
g9953 and b[31] n2198 ; n10209
g9954 and b[32] n2043 ; n10210
g9955 and n10209_not n10210_not ; n10211
g9956 and n10208_not n10211 ; n10212
g9957 and n2051 n4223 ; n10213
g9958 and n10212 n10213_not ; n10214
g9959 and a[23] n10214_not ; n10215
g9960 and a[23] n10215_not ; n10216
g9961 and n10214_not n10215_not ; n10217
g9962 and n10216_not n10217_not ; n10218
g9963 and n10207 n10218_not ; n10219
g9964 and n10207 n10219_not ; n10220
g9965 and n10218_not n10219_not ; n10221
g9966 and n10220_not n10221_not ; n10222
g9967 and n10018_not n10222 ; n10223
g9968 and n10018 n10222_not ; n10224
g9969 and n10223_not n10224_not ; n10225
g9970 and b[36] n1627 ; n10226
g9971 and b[34] n1763 ; n10227
g9972 and b[35] n1622 ; n10228
g9973 and n10227_not n10228_not ; n10229
g9974 and n10226_not n10229 ; n10230
g9975 and n1630 n4922 ; n10231
g9976 and n10230 n10231_not ; n10232
g9977 and a[20] n10232_not ; n10233
g9978 and a[20] n10233_not ; n10234
g9979 and n10232_not n10233_not ; n10235
g9980 and n10234_not n10235_not ; n10236
g9981 and n10225_not n10236_not ; n10237
g9982 and n10225 n10236 ; n10238
g9983 and n10237_not n10238_not ; n10239
g9984 and n10017 n10239_not ; n10240
g9985 and n10017_not n10239 ; n10241
g9986 and n10240_not n10241_not ; n10242
g9987 and b[39] n1302 ; n10243
g9988 and b[37] n1391 ; n10244
g9989 and b[38] n1297 ; n10245
g9990 and n10244_not n10245_not ; n10246
g9991 and n10243_not n10246 ; n10247
g9992 and n1305 n5451 ; n10248
g9993 and n10247 n10248_not ; n10249
g9994 and a[17] n10249_not ; n10250
g9995 and a[17] n10250_not ; n10251
g9996 and n10249_not n10250_not ; n10252
g9997 and n10251_not n10252_not ; n10253
g9998 and n10242 n10253_not ; n10254
g9999 and n10242 n10254_not ; n10255
g10000 and n10253_not n10254_not ; n10256
g10001 and n10255_not n10256_not ; n10257
g10002 and n9877_not n9883_not ; n10258
g10003 and n10257 n10258 ; n10259
g10004 and n10257_not n10258_not ; n10260
g10005 and n10259_not n10260_not ; n10261
g10006 and b[42] n951 ; n10262
g10007 and b[40] n1056 ; n10263
g10008 and b[41] n946 ; n10264
g10009 and n10263_not n10264_not ; n10265
g10010 and n10262_not n10265 ; n10266
g10011 and n954 n6489 ; n10267
g10012 and n10266 n10267_not ; n10268
g10013 and a[14] n10268_not ; n10269
g10014 and a[14] n10269_not ; n10270
g10015 and n10268_not n10269_not ; n10271
g10016 and n10270_not n10271_not ; n10272
g10017 and n10261_not n10272 ; n10273
g10018 and n10261 n10272_not ; n10274
g10019 and n10273_not n10274_not ; n10275
g10020 and n10016_not n10275 ; n10276
g10021 and n10016 n10275_not ; n10277
g10022 and n10276_not n10277_not ; n10278
g10023 and n10015_not n10278 ; n10279
g10024 and n10015_not n10279_not ; n10280
g10025 and n10278 n10279_not ; n10281
g10026 and n10280_not n10281_not ; n10282
g10027 and n9920_not n10282_not ; n10283
g10028 and n9920_not n10283_not ; n10284
g10029 and n10282_not n10283_not ; n10285
g10030 and n10284_not n10285_not ; n10286
g10031 and b[48] n511 ; n10287
g10032 and b[46] n541 ; n10288
g10033 and b[47] n506 ; n10289
g10034 and n10288_not n10289_not ; n10290
g10035 and n10287_not n10290 ; n10291
g10036 and n514 n8009 ; n10292
g10037 and n10291 n10292_not ; n10293
g10038 and a[8] n10293_not ; n10294
g10039 and a[8] n10294_not ; n10295
g10040 and n10293_not n10294_not ; n10296
g10041 and n10295_not n10296_not ; n10297
g10042 and n10286_not n10297_not ; n10298
g10043 and n10286_not n10298_not ; n10299
g10044 and n10297_not n10298_not ; n10300
g10045 and n10299_not n10300_not ; n10301
g10046 and n9934_not n9940_not ; n10302
g10047 and n10301 n10302 ; n10303
g10048 and n10301_not n10302_not ; n10304
g10049 and n10303_not n10304_not ; n10305
g10050 and b[51] n362 ; n10306
g10051 and b[49] n403 ; n10307
g10052 and b[50] n357 ; n10308
g10053 and n10307_not n10308_not ; n10309
g10054 and n10306_not n10309 ; n10310
g10055 and n365 n8976 ; n10311
g10056 and n10310 n10311_not ; n10312
g10057 and a[5] n10312_not ; n10313
g10058 and a[5] n10313_not ; n10314
g10059 and n10312_not n10313_not ; n10315
g10060 and n10314_not n10315_not ; n10316
g10061 and n10305_not n10316 ; n10317
g10062 and n10305 n10316_not ; n10318
g10063 and n10317_not n10318_not ; n10319
g10064 and n9958_not n10319 ; n10320
g10065 and n9958 n10319_not ; n10321
g10066 and n10320_not n10321_not ; n10322
g10067 and n10004_not n10322 ; n10323
g10068 and n10004 n10322_not ; n10324
g10069 and n10323_not n10324_not ; n10325
g10070 and n9986_not n10325 ; n10326
g10071 and n9986 n10325_not ; n10327
g10072 and n10326_not n10327_not ; f[54]
g10073 and n10323_not n10326_not ; n10329
g10074 and n10318_not n10320_not ; n10330
g10075 and b[52] n362 ; n10331
g10076 and b[50] n403 ; n10332
g10077 and b[51] n357 ; n10333
g10078 and n10332_not n10333_not ; n10334
g10079 and n10331_not n10334 ; n10335
g10080 and n365 n9628 ; n10336
g10081 and n10335 n10336_not ; n10337
g10082 and a[5] n10337_not ; n10338
g10083 and a[5] n10338_not ; n10339
g10084 and n10337_not n10338_not ; n10340
g10085 and n10339_not n10340_not ; n10341
g10086 and n10298_not n10304_not ; n10342
g10087 and b[49] n511 ; n10343
g10088 and b[47] n541 ; n10344
g10089 and b[48] n506 ; n10345
g10090 and n10344_not n10345_not ; n10346
g10091 and n10343_not n10346 ; n10347
g10092 and n514 n8625 ; n10348
g10093 and n10347 n10348_not ; n10349
g10094 and a[8] n10349_not ; n10350
g10095 and a[8] n10350_not ; n10351
g10096 and n10349_not n10350_not ; n10352
g10097 and n10351_not n10352_not ; n10353
g10098 and n10279_not n10283_not ; n10354
g10099 and n10274_not n10276_not ; n10355
g10100 and n10176_not n10180_not ; n10356
g10101 and b[16] n5777 ; n10357
g10102 and b[14] n6059 ; n10358
g10103 and b[15] n5772 ; n10359
g10104 and n10358_not n10359_not ; n10360
g10105 and n10357_not n10360 ; n10361
g10106 and n1237 n5780 ; n10362
g10107 and n10361 n10362_not ; n10363
g10108 and a[41] n10363_not ; n10364
g10109 and a[41] n10364_not ; n10365
g10110 and n10363_not n10364_not ; n10366
g10111 and n10365_not n10366_not ; n10367
g10112 and n10162_not n10166_not ; n10368
g10113 and b[13] n6595 ; n10369
g10114 and b[11] n6902 ; n10370
g10115 and b[12] n6590 ; n10371
g10116 and n10370_not n10371_not ; n10372
g10117 and n10369_not n10372 ; n10373
g10118 and n1008 n6598 ; n10374
g10119 and n10373 n10374_not ; n10375
g10120 and a[44] n10375_not ; n10376
g10121 and a[44] n10376_not ; n10377
g10122 and n10375_not n10376_not ; n10378
g10123 and n10377_not n10378_not ; n10379
g10124 and n10154_not n10158_not ; n10380
g10125 and b[10] n7446 ; n10381
g10126 and b[8] n7787 ; n10382
g10127 and b[9] n7441 ; n10383
g10128 and n10382_not n10383_not ; n10384
g10129 and n10381_not n10384 ; n10385
g10130 and n738 n7449 ; n10386
g10131 and n10385 n10386_not ; n10387
g10132 and a[47] n10387_not ; n10388
g10133 and a[47] n10388_not ; n10389
g10134 and n10387_not n10388_not ; n10390
g10135 and n10389_not n10390_not ; n10391
g10136 and n10147_not n10151_not ; n10392
g10137 and b[7] n8362 ; n10393
g10138 and b[5] n8715 ; n10394
g10139 and b[6] n8357 ; n10395
g10140 and n10394_not n10395_not ; n10396
g10141 and n10393_not n10396 ; n10397
g10142 and n484 n8365 ; n10398
g10143 and n10397 n10398_not ; n10399
g10144 and a[50] n10399_not ; n10400
g10145 and a[50] n10400_not ; n10401
g10146 and n10399_not n10400_not ; n10402
g10147 and n10401_not n10402_not ; n10403
g10148 and n9744 n10129 ; n10404
g10149 and n10144_not n10404_not ; n10405
g10150 and b[4] n9339 ; n10406
g10151 and b[2] n9732 ; n10407
g10152 and b[3] n9334 ; n10408
g10153 and n10407_not n10408_not ; n10409
g10154 and n10406_not n10409 ; n10410
g10155 and n346 n9342 ; n10411
g10156 and n10410 n10411_not ; n10412
g10157 and a[53] n10412_not ; n10413
g10158 and a[53] n10413_not ; n10414
g10159 and n10412_not n10413_not ; n10415
g10160 and n10414_not n10415_not ; n10416
g10161 and a[56] n10129_not ; n10417
g10162 and a[54]_not a[55] ; n10418
g10163 and a[54] a[55]_not ; n10419
g10164 and n10418_not n10419_not ; n10420
g10165 and n10128 n10420_not ; n10421
g10166 and b[0] n10421 ; n10422
g10167 and a[55]_not a[56] ; n10423
g10168 and a[55] a[56]_not ; n10424
g10169 and n10423_not n10424_not ; n10425
g10170 and n10128_not n10425 ; n10426
g10171 and b[1] n10426 ; n10427
g10172 and n10422_not n10427_not ; n10428
g10173 and n10128_not n10425_not ; n10429
g10174 and n272_not n10429 ; n10430
g10175 and n10428 n10430_not ; n10431
g10176 and a[56] n10431_not ; n10432
g10177 and a[56] n10432_not ; n10433
g10178 and n10431_not n10432_not ; n10434
g10179 and n10433_not n10434_not ; n10435
g10180 and n10417 n10435_not ; n10436
g10181 and n10417_not n10435 ; n10437
g10182 and n10436_not n10437_not ; n10438
g10183 and n10416 n10438_not ; n10439
g10184 and n10416_not n10438 ; n10440
g10185 and n10439_not n10440_not ; n10441
g10186 and n10405_not n10441 ; n10442
g10187 and n10405 n10441_not ; n10443
g10188 and n10442_not n10443_not ; n10444
g10189 and n10403 n10444_not ; n10445
g10190 and n10403_not n10444 ; n10446
g10191 and n10445_not n10446_not ; n10447
g10192 and n10392_not n10447 ; n10448
g10193 and n10392 n10447_not ; n10449
g10194 and n10448_not n10449_not ; n10450
g10195 and n10391 n10450_not ; n10451
g10196 and n10391_not n10450 ; n10452
g10197 and n10451_not n10452_not ; n10453
g10198 and n10380_not n10453 ; n10454
g10199 and n10380 n10453_not ; n10455
g10200 and n10454_not n10455_not ; n10456
g10201 and n10379 n10456_not ; n10457
g10202 and n10379_not n10456 ; n10458
g10203 and n10457_not n10458_not ; n10459
g10204 and n10368_not n10459 ; n10460
g10205 and n10368 n10459_not ; n10461
g10206 and n10460_not n10461_not ; n10462
g10207 and n10367_not n10462 ; n10463
g10208 and n10462 n10463_not ; n10464
g10209 and n10367_not n10463_not ; n10465
g10210 and n10464_not n10465_not ; n10466
g10211 and n10170_not n10173_not ; n10467
g10212 and n10466 n10467 ; n10468
g10213 and n10466_not n10467_not ; n10469
g10214 and n10468_not n10469_not ; n10470
g10215 and b[19] n5035 ; n10471
g10216 and b[17] n5277 ; n10472
g10217 and b[18] n5030 ; n10473
g10218 and n10472_not n10473_not ; n10474
g10219 and n10471_not n10474 ; n10475
g10220 and n1708 n5038 ; n10476
g10221 and n10475 n10476_not ; n10477
g10222 and a[38] n10477_not ; n10478
g10223 and a[38] n10478_not ; n10479
g10224 and n10477_not n10478_not ; n10480
g10225 and n10479_not n10480_not ; n10481
g10226 and n10470 n10481_not ; n10482
g10227 and n10470_not n10481 ; n10483
g10228 and n10356_not n10483_not ; n10484
g10229 and n10482_not n10484 ; n10485
g10230 and n10356_not n10485_not ; n10486
g10231 and n10482_not n10485_not ; n10487
g10232 and n10483_not n10487 ; n10488
g10233 and n10486_not n10488_not ; n10489
g10234 and b[22] n4287 ; n10490
g10235 and b[20] n4532 ; n10491
g10236 and b[21] n4282 ; n10492
g10237 and n10491_not n10492_not ; n10493
g10238 and n10490_not n10493 ; n10494
g10239 and n2145 n4290 ; n10495
g10240 and n10494 n10495_not ; n10496
g10241 and a[35] n10496_not ; n10497
g10242 and a[35] n10497_not ; n10498
g10243 and n10496_not n10497_not ; n10499
g10244 and n10498_not n10499_not ; n10500
g10245 and n10489_not n10500_not ; n10501
g10246 and n10489_not n10501_not ; n10502
g10247 and n10500_not n10501_not ; n10503
g10248 and n10502_not n10503_not ; n10504
g10249 and n10184_not n10187_not ; n10505
g10250 and n10504 n10505 ; n10506
g10251 and n10504_not n10505_not ; n10507
g10252 and n10506_not n10507_not ; n10508
g10253 and b[25] n3638 ; n10509
g10254 and b[23] n3843 ; n10510
g10255 and b[24] n3633 ; n10511
g10256 and n10510_not n10511_not ; n10512
g10257 and n10509_not n10512 ; n10513
g10258 and n2485 n3641 ; n10514
g10259 and n10513 n10514_not ; n10515
g10260 and a[32] n10515_not ; n10516
g10261 and a[32] n10516_not ; n10517
g10262 and n10515_not n10516_not ; n10518
g10263 and n10517_not n10518_not ; n10519
g10264 and n10508 n10519_not ; n10520
g10265 and n10508 n10520_not ; n10521
g10266 and n10519_not n10520_not ; n10522
g10267 and n10521_not n10522_not ; n10523
g10268 and n10190_not n10193_not ; n10524
g10269 and n10523 n10524 ; n10525
g10270 and n10523_not n10524_not ; n10526
g10271 and n10525_not n10526_not ; n10527
g10272 and b[28] n3050 ; n10528
g10273 and b[26] n3243 ; n10529
g10274 and b[27] n3045 ; n10530
g10275 and n10529_not n10530_not ; n10531
g10276 and n10528_not n10531 ; n10532
g10277 and n3053 n3189 ; n10533
g10278 and n10532 n10533_not ; n10534
g10279 and a[29] n10534_not ; n10535
g10280 and a[29] n10535_not ; n10536
g10281 and n10534_not n10535_not ; n10537
g10282 and n10536_not n10537_not ; n10538
g10283 and n10527 n10538_not ; n10539
g10284 and n10527 n10539_not ; n10540
g10285 and n10538_not n10539_not ; n10541
g10286 and n10540_not n10541_not ; n10542
g10287 and n10196_not n10199_not ; n10543
g10288 and n10542 n10543 ; n10544
g10289 and n10542_not n10543_not ; n10545
g10290 and n10544_not n10545_not ; n10546
g10291 and b[31] n2539 ; n10547
g10292 and b[29] n2685 ; n10548
g10293 and b[30] n2534 ; n10549
g10294 and n10548_not n10549_not ; n10550
g10295 and n10547_not n10550 ; n10551
g10296 and n2542 n3796 ; n10552
g10297 and n10551 n10552_not ; n10553
g10298 and a[26] n10553_not ; n10554
g10299 and a[26] n10554_not ; n10555
g10300 and n10553_not n10554_not ; n10556
g10301 and n10555_not n10556_not ; n10557
g10302 and n10546 n10557_not ; n10558
g10303 and n10546 n10558_not ; n10559
g10304 and n10557_not n10558_not ; n10560
g10305 and n10559_not n10560_not ; n10561
g10306 and n10202_not n10205_not ; n10562
g10307 and n10561 n10562 ; n10563
g10308 and n10561_not n10562_not ; n10564
g10309 and n10563_not n10564_not ; n10565
g10310 and b[34] n2048 ; n10566
g10311 and b[32] n2198 ; n10567
g10312 and b[33] n2043 ; n10568
g10313 and n10567_not n10568_not ; n10569
g10314 and n10566_not n10569 ; n10570
g10315 and n2051 n4466 ; n10571
g10316 and n10570 n10571_not ; n10572
g10317 and a[23] n10572_not ; n10573
g10318 and a[23] n10573_not ; n10574
g10319 and n10572_not n10573_not ; n10575
g10320 and n10574_not n10575_not ; n10576
g10321 and n10565 n10576_not ; n10577
g10322 and n10565 n10577_not ; n10578
g10323 and n10576_not n10577_not ; n10579
g10324 and n10578_not n10579_not ; n10580
g10325 and n10018_not n10222_not ; n10581
g10326 and n10219_not n10581_not ; n10582
g10327 and n10580 n10582 ; n10583
g10328 and n10580_not n10582_not ; n10584
g10329 and n10583_not n10584_not ; n10585
g10330 and b[37] n1627 ; n10586
g10331 and b[35] n1763 ; n10587
g10332 and b[36] n1622 ; n10588
g10333 and n10587_not n10588_not ; n10589
g10334 and n10586_not n10589 ; n10590
g10335 and n1630 n5181 ; n10591
g10336 and n10590 n10591_not ; n10592
g10337 and a[20] n10592_not ; n10593
g10338 and a[20] n10593_not ; n10594
g10339 and n10592_not n10593_not ; n10595
g10340 and n10594_not n10595_not ; n10596
g10341 and n10585 n10596_not ; n10597
g10342 and n10585 n10597_not ; n10598
g10343 and n10596_not n10597_not ; n10599
g10344 and n10598_not n10599_not ; n10600
g10345 and n10237_not n10241_not ; n10601
g10346 and n10600 n10601 ; n10602
g10347 and n10600_not n10601_not ; n10603
g10348 and n10602_not n10603_not ; n10604
g10349 and b[40] n1302 ; n10605
g10350 and b[38] n1391 ; n10606
g10351 and b[39] n1297 ; n10607
g10352 and n10606_not n10607_not ; n10608
g10353 and n10605_not n10608 ; n10609
g10354 and n1305 n5955 ; n10610
g10355 and n10609 n10610_not ; n10611
g10356 and a[17] n10611_not ; n10612
g10357 and a[17] n10612_not ; n10613
g10358 and n10611_not n10612_not ; n10614
g10359 and n10613_not n10614_not ; n10615
g10360 and n10604 n10615_not ; n10616
g10361 and n10604 n10616_not ; n10617
g10362 and n10615_not n10616_not ; n10618
g10363 and n10617_not n10618_not ; n10619
g10364 and n10254_not n10260_not ; n10620
g10365 and n10619 n10620 ; n10621
g10366 and n10619_not n10620_not ; n10622
g10367 and n10621_not n10622_not ; n10623
g10368 and b[43] n951 ; n10624
g10369 and b[41] n1056 ; n10625
g10370 and b[42] n946 ; n10626
g10371 and n10625_not n10626_not ; n10627
g10372 and n10624_not n10627 ; n10628
g10373 and n954 n6515 ; n10629
g10374 and n10628 n10629_not ; n10630
g10375 and a[14] n10630_not ; n10631
g10376 and a[14] n10631_not ; n10632
g10377 and n10630_not n10631_not ; n10633
g10378 and n10632_not n10633_not ; n10634
g10379 and n10623 n10634_not ; n10635
g10380 and n10623_not n10634 ; n10636
g10381 and n10355_not n10636_not ; n10637
g10382 and n10635_not n10637 ; n10638
g10383 and n10355_not n10638_not ; n10639
g10384 and n10635_not n10638_not ; n10640
g10385 and n10636_not n10640 ; n10641
g10386 and n10639_not n10641_not ; n10642
g10387 and b[46] n700 ; n10643
g10388 and b[44] n767 ; n10644
g10389 and b[45] n695 ; n10645
g10390 and n10644_not n10645_not ; n10646
g10391 and n10643_not n10646 ; n10647
g10392 and n703 n7677 ; n10648
g10393 and n10647 n10648_not ; n10649
g10394 and a[11] n10649_not ; n10650
g10395 and a[11] n10650_not ; n10651
g10396 and n10649_not n10650_not ; n10652
g10397 and n10651_not n10652_not ; n10653
g10398 and n10642 n10653 ; n10654
g10399 and n10642_not n10653_not ; n10655
g10400 and n10654_not n10655_not ; n10656
g10401 and n10354_not n10656 ; n10657
g10402 and n10354 n10656_not ; n10658
g10403 and n10657_not n10658_not ; n10659
g10404 and n10353 n10659_not ; n10660
g10405 and n10353_not n10659 ; n10661
g10406 and n10660_not n10661_not ; n10662
g10407 and n10342_not n10662 ; n10663
g10408 and n10342 n10662_not ; n10664
g10409 and n10663_not n10664_not ; n10665
g10410 and n10341_not n10665 ; n10666
g10411 and n10665 n10666_not ; n10667
g10412 and n10341_not n10666_not ; n10668
g10413 and n10667_not n10668_not ; n10669
g10414 and n10330_not n10669 ; n10670
g10415 and n10330 n10669_not ; n10671
g10416 and n10670_not n10671_not ; n10672
g10417 and b[55] n266 ; n10673
g10418 and b[53] n284 ; n10674
g10419 and b[54] n261 ; n10675
g10420 and n10674_not n10675_not ; n10676
g10421 and n10673_not n10676 ; n10677
g10422 and n9994_not n9996_not ; n10678
g10423 and b[54]_not b[55]_not ; n10679
g10424 and b[54] b[55] ; n10680
g10425 and n10679_not n10680_not ; n10681
g10426 and n10678_not n10681 ; n10682
g10427 and n10678 n10681_not ; n10683
g10428 and n10682_not n10683_not ; n10684
g10429 and n269 n10684 ; n10685
g10430 and n10677 n10685_not ; n10686
g10431 and a[2] n10686_not ; n10687
g10432 and a[2] n10687_not ; n10688
g10433 and n10686_not n10687_not ; n10689
g10434 and n10688_not n10689_not ; n10690
g10435 and n10672_not n10690_not ; n10691
g10436 and n10672 n10690 ; n10692
g10437 and n10691_not n10692_not ; n10693
g10438 and n10329_not n10693 ; n10694
g10439 and n10329 n10693_not ; n10695
g10440 and n10694_not n10695_not ; f[55]
g10441 and b[56] n266 ; n10697
g10442 and b[54] n284 ; n10698
g10443 and b[55] n261 ; n10699
g10444 and n10698_not n10699_not ; n10700
g10445 and n10697_not n10700 ; n10701
g10446 and n10680_not n10682_not ; n10702
g10447 and b[55]_not b[56]_not ; n10703
g10448 and b[55] b[56] ; n10704
g10449 and n10703_not n10704_not ; n10705
g10450 and n10702_not n10705 ; n10706
g10451 and n10702 n10705_not ; n10707
g10452 and n10706_not n10707_not ; n10708
g10453 and n269 n10708 ; n10709
g10454 and n10701 n10709_not ; n10710
g10455 and a[2] n10710_not ; n10711
g10456 and a[2] n10711_not ; n10712
g10457 and n10710_not n10711_not ; n10713
g10458 and n10712_not n10713_not ; n10714
g10459 and n10330_not n10669_not ; n10715
g10460 and n10666_not n10715_not ; n10716
g10461 and n10661_not n10663_not ; n10717
g10462 and b[50] n511 ; n10718
g10463 and b[48] n541 ; n10719
g10464 and b[49] n506 ; n10720
g10465 and n10719_not n10720_not ; n10721
g10466 and n10718_not n10721 ; n10722
g10467 and n514 n8949 ; n10723
g10468 and n10722 n10723_not ; n10724
g10469 and a[8] n10724_not ; n10725
g10470 and a[8] n10725_not ; n10726
g10471 and n10724_not n10725_not ; n10727
g10472 and n10726_not n10727_not ; n10728
g10473 and n10655_not n10657_not ; n10729
g10474 and b[35] n2048 ; n10730
g10475 and b[33] n2198 ; n10731
g10476 and b[34] n2043 ; n10732
g10477 and n10731_not n10732_not ; n10733
g10478 and n10730_not n10733 ; n10734
g10479 and n2051 n4696 ; n10735
g10480 and n10734 n10735_not ; n10736
g10481 and a[23] n10736_not ; n10737
g10482 and a[23] n10737_not ; n10738
g10483 and n10736_not n10737_not ; n10739
g10484 and n10738_not n10739_not ; n10740
g10485 and n10558_not n10564_not ; n10741
g10486 and b[32] n2539 ; n10742
g10487 and b[30] n2685 ; n10743
g10488 and b[31] n2534 ; n10744
g10489 and n10743_not n10744_not ; n10745
g10490 and n10742_not n10745 ; n10746
g10491 and n2542 n4013 ; n10747
g10492 and n10746 n10747_not ; n10748
g10493 and a[26] n10748_not ; n10749
g10494 and a[26] n10749_not ; n10750
g10495 and n10748_not n10749_not ; n10751
g10496 and n10750_not n10751_not ; n10752
g10497 and n10539_not n10545_not ; n10753
g10498 and n10520_not n10526_not ; n10754
g10499 and n10501_not n10507_not ; n10755
g10500 and n10463_not n10469_not ; n10756
g10501 and b[17] n5777 ; n10757
g10502 and b[15] n6059 ; n10758
g10503 and b[16] n5772 ; n10759
g10504 and n10758_not n10759_not ; n10760
g10505 and n10757_not n10760 ; n10761
g10506 and n1356 n5780 ; n10762
g10507 and n10761 n10762_not ; n10763
g10508 and a[41] n10763_not ; n10764
g10509 and a[41] n10764_not ; n10765
g10510 and n10763_not n10764_not ; n10766
g10511 and n10765_not n10766_not ; n10767
g10512 and n10458_not n10460_not ; n10768
g10513 and b[14] n6595 ; n10769
g10514 and b[12] n6902 ; n10770
g10515 and b[13] n6590 ; n10771
g10516 and n10770_not n10771_not ; n10772
g10517 and n10769_not n10772 ; n10773
g10518 and n1034 n6598 ; n10774
g10519 and n10773 n10774_not ; n10775
g10520 and a[44] n10775_not ; n10776
g10521 and a[44] n10776_not ; n10777
g10522 and n10775_not n10776_not ; n10778
g10523 and n10777_not n10778_not ; n10779
g10524 and n10452_not n10454_not ; n10780
g10525 and b[11] n7446 ; n10781
g10526 and b[9] n7787 ; n10782
g10527 and b[10] n7441 ; n10783
g10528 and n10782_not n10783_not ; n10784
g10529 and n10781_not n10784 ; n10785
g10530 and n818 n7449 ; n10786
g10531 and n10785 n10786_not ; n10787
g10532 and a[47] n10787_not ; n10788
g10533 and a[47] n10788_not ; n10789
g10534 and n10787_not n10788_not ; n10790
g10535 and n10789_not n10790_not ; n10791
g10536 and n10446_not n10448_not ; n10792
g10537 and n10440_not n10442_not ; n10793
g10538 and b[2] n10426 ; n10794
g10539 and n10128 n10425_not ; n10795
g10540 and n10420 n10795 ; n10796
g10541 and b[0] n10796 ; n10797
g10542 and b[1] n10421 ; n10798
g10543 and n10797_not n10798_not ; n10799
g10544 and n10794_not n10799 ; n10800
g10545 and n296 n10429 ; n10801
g10546 and n10800 n10801_not ; n10802
g10547 and a[56] n10802_not ; n10803
g10548 and a[56] n10803_not ; n10804
g10549 and n10802_not n10803_not ; n10805
g10550 and n10804_not n10805_not ; n10806
g10551 and n10436_not n10806 ; n10807
g10552 and n10436 n10806_not ; n10808
g10553 and n10807_not n10808_not ; n10809
g10554 and b[5] n9339 ; n10810
g10555 and b[3] n9732 ; n10811
g10556 and b[4] n9334 ; n10812
g10557 and n10811_not n10812_not ; n10813
g10558 and n10810_not n10813 ; n10814
g10559 and n394 n9342 ; n10815
g10560 and n10814 n10815_not ; n10816
g10561 and a[53] n10816_not ; n10817
g10562 and a[53] n10817_not ; n10818
g10563 and n10816_not n10817_not ; n10819
g10564 and n10818_not n10819_not ; n10820
g10565 and n10809 n10820_not ; n10821
g10566 and n10809_not n10820 ; n10822
g10567 and n10793_not n10822_not ; n10823
g10568 and n10821_not n10823 ; n10824
g10569 and n10793_not n10824_not ; n10825
g10570 and n10821_not n10824_not ; n10826
g10571 and n10822_not n10826 ; n10827
g10572 and n10825_not n10827_not ; n10828
g10573 and b[8] n8362 ; n10829
g10574 and b[6] n8715 ; n10830
g10575 and b[7] n8357 ; n10831
g10576 and n10830_not n10831_not ; n10832
g10577 and n10829_not n10832 ; n10833
g10578 and n585 n8365 ; n10834
g10579 and n10833 n10834_not ; n10835
g10580 and a[50] n10835_not ; n10836
g10581 and a[50] n10836_not ; n10837
g10582 and n10835_not n10836_not ; n10838
g10583 and n10837_not n10838_not ; n10839
g10584 and n10828 n10839 ; n10840
g10585 and n10828_not n10839_not ; n10841
g10586 and n10840_not n10841_not ; n10842
g10587 and n10792_not n10842 ; n10843
g10588 and n10792 n10842_not ; n10844
g10589 and n10843_not n10844_not ; n10845
g10590 and n10791 n10845_not ; n10846
g10591 and n10791_not n10845 ; n10847
g10592 and n10846_not n10847_not ; n10848
g10593 and n10780_not n10848 ; n10849
g10594 and n10780 n10848_not ; n10850
g10595 and n10849_not n10850_not ; n10851
g10596 and n10779_not n10851 ; n10852
g10597 and n10851 n10852_not ; n10853
g10598 and n10779_not n10852_not ; n10854
g10599 and n10853_not n10854_not ; n10855
g10600 and n10768_not n10855_not ; n10856
g10601 and n10768 n10855 ; n10857
g10602 and n10856_not n10857_not ; n10858
g10603 and n10767_not n10858 ; n10859
g10604 and n10767_not n10859_not ; n10860
g10605 and n10858 n10859_not ; n10861
g10606 and n10860_not n10861_not ; n10862
g10607 and n10756_not n10862_not ; n10863
g10608 and n10756_not n10863_not ; n10864
g10609 and n10862_not n10863_not ; n10865
g10610 and n10864_not n10865_not ; n10866
g10611 and b[20] n5035 ; n10867
g10612 and b[18] n5277 ; n10868
g10613 and b[19] n5030 ; n10869
g10614 and n10868_not n10869_not ; n10870
g10615 and n10867_not n10870 ; n10871
g10616 and n1846 n5038 ; n10872
g10617 and n10871 n10872_not ; n10873
g10618 and a[38] n10873_not ; n10874
g10619 and a[38] n10874_not ; n10875
g10620 and n10873_not n10874_not ; n10876
g10621 and n10875_not n10876_not ; n10877
g10622 and n10866_not n10877_not ; n10878
g10623 and n10866_not n10878_not ; n10879
g10624 and n10877_not n10878_not ; n10880
g10625 and n10879_not n10880_not ; n10881
g10626 and n10487_not n10881 ; n10882
g10627 and n10487 n10881_not ; n10883
g10628 and n10882_not n10883_not ; n10884
g10629 and b[23] n4287 ; n10885
g10630 and b[21] n4532 ; n10886
g10631 and b[22] n4282 ; n10887
g10632 and n10886_not n10887_not ; n10888
g10633 and n10885_not n10888 ; n10889
g10634 and n2300 n4290 ; n10890
g10635 and n10889 n10890_not ; n10891
g10636 and a[35] n10891_not ; n10892
g10637 and a[35] n10892_not ; n10893
g10638 and n10891_not n10892_not ; n10894
g10639 and n10893_not n10894_not ; n10895
g10640 and n10884_not n10895_not ; n10896
g10641 and n10884 n10895 ; n10897
g10642 and n10896_not n10897_not ; n10898
g10643 and n10755 n10898_not ; n10899
g10644 and n10755_not n10898 ; n10900
g10645 and n10899_not n10900_not ; n10901
g10646 and b[26] n3638 ; n10902
g10647 and b[24] n3843 ; n10903
g10648 and b[25] n3633 ; n10904
g10649 and n10903_not n10904_not ; n10905
g10650 and n10902_not n10905 ; n10906
g10651 and n2813 n3641 ; n10907
g10652 and n10906 n10907_not ; n10908
g10653 and a[32] n10908_not ; n10909
g10654 and a[32] n10909_not ; n10910
g10655 and n10908_not n10909_not ; n10911
g10656 and n10910_not n10911_not ; n10912
g10657 and n10901 n10912_not ; n10913
g10658 and n10901_not n10912 ; n10914
g10659 and n10754_not n10914_not ; n10915
g10660 and n10913_not n10915 ; n10916
g10661 and n10754_not n10916_not ; n10917
g10662 and n10913_not n10916_not ; n10918
g10663 and n10914_not n10918 ; n10919
g10664 and n10917_not n10919_not ; n10920
g10665 and b[29] n3050 ; n10921
g10666 and b[27] n3243 ; n10922
g10667 and b[28] n3045 ; n10923
g10668 and n10922_not n10923_not ; n10924
g10669 and n10921_not n10924 ; n10925
g10670 and n3053 n3383 ; n10926
g10671 and n10925 n10926_not ; n10927
g10672 and a[29] n10927_not ; n10928
g10673 and a[29] n10928_not ; n10929
g10674 and n10927_not n10928_not ; n10930
g10675 and n10929_not n10930_not ; n10931
g10676 and n10920 n10931 ; n10932
g10677 and n10920_not n10931_not ; n10933
g10678 and n10932_not n10933_not ; n10934
g10679 and n10753_not n10934 ; n10935
g10680 and n10753 n10934_not ; n10936
g10681 and n10935_not n10936_not ; n10937
g10682 and n10752 n10937_not ; n10938
g10683 and n10752_not n10937 ; n10939
g10684 and n10938_not n10939_not ; n10940
g10685 and n10741_not n10940 ; n10941
g10686 and n10741 n10940_not ; n10942
g10687 and n10941_not n10942_not ; n10943
g10688 and n10740_not n10943 ; n10944
g10689 and n10943 n10944_not ; n10945
g10690 and n10740_not n10944_not ; n10946
g10691 and n10945_not n10946_not ; n10947
g10692 and n10577_not n10584_not ; n10948
g10693 and n10947 n10948 ; n10949
g10694 and n10947_not n10948_not ; n10950
g10695 and n10949_not n10950_not ; n10951
g10696 and b[38] n1627 ; n10952
g10697 and b[36] n1763 ; n10953
g10698 and b[37] n1622 ; n10954
g10699 and n10953_not n10954_not ; n10955
g10700 and n10952_not n10955 ; n10956
g10701 and n1630 n5205 ; n10957
g10702 and n10956 n10957_not ; n10958
g10703 and a[20] n10958_not ; n10959
g10704 and a[20] n10959_not ; n10960
g10705 and n10958_not n10959_not ; n10961
g10706 and n10960_not n10961_not ; n10962
g10707 and n10951 n10962_not ; n10963
g10708 and n10951 n10963_not ; n10964
g10709 and n10962_not n10963_not ; n10965
g10710 and n10964_not n10965_not ; n10966
g10711 and n10597_not n10603_not ; n10967
g10712 and n10966 n10967 ; n10968
g10713 and n10966_not n10967_not ; n10969
g10714 and n10968_not n10969_not ; n10970
g10715 and b[41] n1302 ; n10971
g10716 and b[39] n1391 ; n10972
g10717 and b[40] n1297 ; n10973
g10718 and n10972_not n10973_not ; n10974
g10719 and n10971_not n10974 ; n10975
g10720 and n1305 n6219 ; n10976
g10721 and n10975 n10976_not ; n10977
g10722 and a[17] n10977_not ; n10978
g10723 and a[17] n10978_not ; n10979
g10724 and n10977_not n10978_not ; n10980
g10725 and n10979_not n10980_not ; n10981
g10726 and n10970 n10981_not ; n10982
g10727 and n10970 n10982_not ; n10983
g10728 and n10981_not n10982_not ; n10984
g10729 and n10983_not n10984_not ; n10985
g10730 and n10616_not n10622_not ; n10986
g10731 and n10985 n10986 ; n10987
g10732 and n10985_not n10986_not ; n10988
g10733 and n10987_not n10988_not ; n10989
g10734 and b[44] n951 ; n10990
g10735 and b[42] n1056 ; n10991
g10736 and b[43] n946 ; n10992
g10737 and n10991_not n10992_not ; n10993
g10738 and n10990_not n10993 ; n10994
g10739 and n954 n7072 ; n10995
g10740 and n10994 n10995_not ; n10996
g10741 and a[14] n10996_not ; n10997
g10742 and a[14] n10997_not ; n10998
g10743 and n10996_not n10997_not ; n10999
g10744 and n10998_not n10999_not ; n11000
g10745 and n10989 n11000_not ; n11001
g10746 and n10989_not n11000 ; n11002
g10747 and n10640_not n11002_not ; n11003
g10748 and n11001_not n11003 ; n11004
g10749 and n10640_not n11004_not ; n11005
g10750 and n11001_not n11004_not ; n11006
g10751 and n11002_not n11006 ; n11007
g10752 and n11005_not n11007_not ; n11008
g10753 and b[47] n700 ; n11009
g10754 and b[45] n767 ; n11010
g10755 and b[46] n695 ; n11011
g10756 and n11010_not n11011_not ; n11012
g10757 and n11009_not n11012 ; n11013
g10758 and n703 n7703 ; n11014
g10759 and n11013 n11014_not ; n11015
g10760 and a[11] n11015_not ; n11016
g10761 and a[11] n11016_not ; n11017
g10762 and n11015_not n11016_not ; n11018
g10763 and n11017_not n11018_not ; n11019
g10764 and n11008_not n11019_not ; n11020
g10765 and n11008_not n11020_not ; n11021
g10766 and n11019_not n11020_not ; n11022
g10767 and n11021_not n11022_not ; n11023
g10768 and n10729_not n11023_not ; n11024
g10769 and n10729 n11023 ; n11025
g10770 and n11024_not n11025_not ; n11026
g10771 and n10728_not n11026 ; n11027
g10772 and n10728_not n11027_not ; n11028
g10773 and n11026 n11027_not ; n11029
g10774 and n11028_not n11029_not ; n11030
g10775 and n10717_not n11030_not ; n11031
g10776 and n10717_not n11031_not ; n11032
g10777 and n11030_not n11031_not ; n11033
g10778 and n11032_not n11033_not ; n11034
g10779 and b[53] n362 ; n11035
g10780 and b[51] n403 ; n11036
g10781 and b[52] n357 ; n11037
g10782 and n11036_not n11037_not ; n11038
g10783 and n11035_not n11038 ; n11039
g10784 and n365 n9972 ; n11040
g10785 and n11039 n11040_not ; n11041
g10786 and a[5] n11041_not ; n11042
g10787 and a[5] n11042_not ; n11043
g10788 and n11041_not n11042_not ; n11044
g10789 and n11043_not n11044_not ; n11045
g10790 and n11034 n11045 ; n11046
g10791 and n11034_not n11045_not ; n11047
g10792 and n11046_not n11047_not ; n11048
g10793 and n10716_not n11048 ; n11049
g10794 and n10716 n11048_not ; n11050
g10795 and n11049_not n11050_not ; n11051
g10796 and n10714_not n11051 ; n11052
g10797 and n11051 n11052_not ; n11053
g10798 and n10714_not n11052_not ; n11054
g10799 and n11053_not n11054_not ; n11055
g10800 and n10691_not n10694_not ; n11056
g10801 and n11055_not n11056_not ; n11057
g10802 and n11055 n11056 ; n11058
g10803 and n11057_not n11058_not ; f[56]
g10804 and n11047_not n11049_not ; n11060
g10805 and b[54] n362 ; n11061
g10806 and b[52] n403 ; n11062
g10807 and b[53] n357 ; n11063
g10808 and n11062_not n11063_not ; n11064
g10809 and n11061_not n11064 ; n11065
g10810 and n365 n9998 ; n11066
g10811 and n11065 n11066_not ; n11067
g10812 and a[5] n11067_not ; n11068
g10813 and a[5] n11068_not ; n11069
g10814 and n11067_not n11068_not ; n11070
g10815 and n11069_not n11070_not ; n11071
g10816 and n11027_not n11031_not ; n11072
g10817 and b[51] n511 ; n11073
g10818 and b[49] n541 ; n11074
g10819 and b[50] n506 ; n11075
g10820 and n11074_not n11075_not ; n11076
g10821 and n11073_not n11076 ; n11077
g10822 and n514 n8976 ; n11078
g10823 and n11077 n11078_not ; n11079
g10824 and a[8] n11079_not ; n11080
g10825 and a[8] n11080_not ; n11081
g10826 and n11079_not n11080_not ; n11082
g10827 and n11081_not n11082_not ; n11083
g10828 and n11020_not n11024_not ; n11084
g10829 and b[48] n700 ; n11085
g10830 and b[46] n767 ; n11086
g10831 and b[47] n695 ; n11087
g10832 and n11086_not n11087_not ; n11088
g10833 and n11085_not n11088 ; n11089
g10834 and n703 n8009 ; n11090
g10835 and n11089 n11090_not ; n11091
g10836 and a[11] n11091_not ; n11092
g10837 and a[11] n11092_not ; n11093
g10838 and n11091_not n11092_not ; n11094
g10839 and n11093_not n11094_not ; n11095
g10840 and b[45] n951 ; n11096
g10841 and b[43] n1056 ; n11097
g10842 and b[44] n946 ; n11098
g10843 and n11097_not n11098_not ; n11099
g10844 and n11096_not n11099 ; n11100
g10845 and n954 n7361 ; n11101
g10846 and n11100 n11101_not ; n11102
g10847 and a[14] n11102_not ; n11103
g10848 and a[14] n11103_not ; n11104
g10849 and n11102_not n11103_not ; n11105
g10850 and n11104_not n11105_not ; n11106
g10851 and n10982_not n10988_not ; n11107
g10852 and n10944_not n10950_not ; n11108
g10853 and n10939_not n10941_not ; n11109
g10854 and n10933_not n10935_not ; n11110
g10855 and b[30] n3050 ; n11111
g10856 and b[28] n3243 ; n11112
g10857 and b[29] n3045 ; n11113
g10858 and n11112_not n11113_not ; n11114
g10859 and n11111_not n11114 ; n11115
g10860 and n3053 n3577 ; n11116
g10861 and n11115 n11116_not ; n11117
g10862 and a[29] n11117_not ; n11118
g10863 and a[29] n11118_not ; n11119
g10864 and n11117_not n11118_not ; n11120
g10865 and n11119_not n11120_not ; n11121
g10866 and n10487_not n10881_not ; n11122
g10867 and n10878_not n11122_not ; n11123
g10868 and b[21] n5035 ; n11124
g10869 and b[19] n5277 ; n11125
g10870 and b[20] n5030 ; n11126
g10871 and n11125_not n11126_not ; n11127
g10872 and n11124_not n11127 ; n11128
g10873 and n1984 n5038 ; n11129
g10874 and n11128 n11129_not ; n11130
g10875 and a[38] n11130_not ; n11131
g10876 and a[38] n11131_not ; n11132
g10877 and n11130_not n11131_not ; n11133
g10878 and n11132_not n11133_not ; n11134
g10879 and n10859_not n10863_not ; n11135
g10880 and b[18] n5777 ; n11136
g10881 and b[16] n6059 ; n11137
g10882 and b[17] n5772 ; n11138
g10883 and n11137_not n11138_not ; n11139
g10884 and n11136_not n11139 ; n11140
g10885 and n1566 n5780 ; n11141
g10886 and n11140 n11141_not ; n11142
g10887 and a[41] n11142_not ; n11143
g10888 and a[41] n11143_not ; n11144
g10889 and n11142_not n11143_not ; n11145
g10890 and n11144_not n11145_not ; n11146
g10891 and n10852_not n10856_not ; n11147
g10892 and b[15] n6595 ; n11148
g10893 and b[13] n6902 ; n11149
g10894 and b[14] n6590 ; n11150
g10895 and n11149_not n11150_not ; n11151
g10896 and n11148_not n11151 ; n11152
g10897 and n1131 n6598 ; n11153
g10898 and n11152 n11153_not ; n11154
g10899 and a[44] n11154_not ; n11155
g10900 and a[44] n11155_not ; n11156
g10901 and n11154_not n11155_not ; n11157
g10902 and n11156_not n11157_not ; n11158
g10903 and n10847_not n10849_not ; n11159
g10904 and b[12] n7446 ; n11160
g10905 and b[10] n7787 ; n11161
g10906 and b[11] n7441 ; n11162
g10907 and n11161_not n11162_not ; n11163
g10908 and n11160_not n11163 ; n11164
g10909 and n842 n7449 ; n11165
g10910 and n11164 n11165_not ; n11166
g10911 and a[47] n11166_not ; n11167
g10912 and a[47] n11167_not ; n11168
g10913 and n11166_not n11167_not ; n11169
g10914 and n11168_not n11169_not ; n11170
g10915 and n10841_not n10843_not ; n11171
g10916 and b[6] n9339 ; n11172
g10917 and b[4] n9732 ; n11173
g10918 and b[5] n9334 ; n11174
g10919 and n11173_not n11174_not ; n11175
g10920 and n11172_not n11175 ; n11176
g10921 and n459 n9342 ; n11177
g10922 and n11176 n11177_not ; n11178
g10923 and a[53] n11178_not ; n11179
g10924 and a[53] n11179_not ; n11180
g10925 and n11178_not n11179_not ; n11181
g10926 and n11180_not n11181_not ; n11182
g10927 and a[56] a[57]_not ; n11183
g10928 and a[56]_not a[57] ; n11184
g10929 and n11183_not n11184_not ; n11185
g10930 and b[0] n11185_not ; n11186
g10931 and n10808_not n11186 ; n11187
g10932 and n10808 n11186_not ; n11188
g10933 and n11187_not n11188_not ; n11189
g10934 and b[3] n10426 ; n11190
g10935 and b[1] n10796 ; n11191
g10936 and b[2] n10421 ; n11192
g10937 and n11191_not n11192_not ; n11193
g10938 and n11190_not n11193 ; n11194
g10939 and n318 n10429 ; n11195
g10940 and n11194 n11195_not ; n11196
g10941 and a[56] n11196_not ; n11197
g10942 and a[56] n11197_not ; n11198
g10943 and n11196_not n11197_not ; n11199
g10944 and n11198_not n11199_not ; n11200
g10945 and n11189_not n11200_not ; n11201
g10946 and n11189 n11200 ; n11202
g10947 and n11201_not n11202_not ; n11203
g10948 and n11182_not n11203 ; n11204
g10949 and n11203 n11204_not ; n11205
g10950 and n11182_not n11204_not ; n11206
g10951 and n11205_not n11206_not ; n11207
g10952 and n10826_not n11207 ; n11208
g10953 and n10826 n11207_not ; n11209
g10954 and n11208_not n11209_not ; n11210
g10955 and b[9] n8362 ; n11211
g10956 and b[7] n8715 ; n11212
g10957 and b[8] n8357 ; n11213
g10958 and n11212_not n11213_not ; n11214
g10959 and n11211_not n11214 ; n11215
g10960 and n651 n8365 ; n11216
g10961 and n11215 n11216_not ; n11217
g10962 and a[50] n11217_not ; n11218
g10963 and a[50] n11218_not ; n11219
g10964 and n11217_not n11218_not ; n11220
g10965 and n11219_not n11220_not ; n11221
g10966 and n11210_not n11221_not ; n11222
g10967 and n11210 n11221 ; n11223
g10968 and n11222_not n11223_not ; n11224
g10969 and n11171_not n11224 ; n11225
g10970 and n11171 n11224_not ; n11226
g10971 and n11225_not n11226_not ; n11227
g10972 and n11170 n11227_not ; n11228
g10973 and n11170_not n11227 ; n11229
g10974 and n11228_not n11229_not ; n11230
g10975 and n11159_not n11230 ; n11231
g10976 and n11159 n11230_not ; n11232
g10977 and n11231_not n11232_not ; n11233
g10978 and n11158_not n11233 ; n11234
g10979 and n11158 n11233_not ; n11235
g10980 and n11234_not n11235_not ; n11236
g10981 and n11147_not n11236 ; n11237
g10982 and n11147 n11236_not ; n11238
g10983 and n11237_not n11238_not ; n11239
g10984 and n11146_not n11239 ; n11240
g10985 and n11146_not n11240_not ; n11241
g10986 and n11239 n11240_not ; n11242
g10987 and n11241_not n11242_not ; n11243
g10988 and n11135_not n11243_not ; n11244
g10989 and n11135 n11242_not ; n11245
g10990 and n11241_not n11245 ; n11246
g10991 and n11244_not n11246_not ; n11247
g10992 and n11134_not n11247 ; n11248
g10993 and n11134 n11247_not ; n11249
g10994 and n11248_not n11249_not ; n11250
g10995 and n11123_not n11250 ; n11251
g10996 and n11123 n11250_not ; n11252
g10997 and n11251_not n11252_not ; n11253
g10998 and b[24] n4287 ; n11254
g10999 and b[22] n4532 ; n11255
g11000 and b[23] n4282 ; n11256
g11001 and n11255_not n11256_not ; n11257
g11002 and n11254_not n11257 ; n11258
g11003 and n2458 n4290 ; n11259
g11004 and n11258 n11259_not ; n11260
g11005 and a[35] n11260_not ; n11261
g11006 and a[35] n11261_not ; n11262
g11007 and n11260_not n11261_not ; n11263
g11008 and n11262_not n11263_not ; n11264
g11009 and n11253 n11264_not ; n11265
g11010 and n11253 n11265_not ; n11266
g11011 and n11264_not n11265_not ; n11267
g11012 and n11266_not n11267_not ; n11268
g11013 and n10896_not n10900_not ; n11269
g11014 and n11268 n11269 ; n11270
g11015 and n11268_not n11269_not ; n11271
g11016 and n11270_not n11271_not ; n11272
g11017 and b[27] n3638 ; n11273
g11018 and b[25] n3843 ; n11274
g11019 and b[26] n3633 ; n11275
g11020 and n11274_not n11275_not ; n11276
g11021 and n11273_not n11276 ; n11277
g11022 and n2990 n3641 ; n11278
g11023 and n11277 n11278_not ; n11279
g11024 and a[32] n11279_not ; n11280
g11025 and a[32] n11280_not ; n11281
g11026 and n11279_not n11280_not ; n11282
g11027 and n11281_not n11282_not ; n11283
g11028 and n11272_not n11283 ; n11284
g11029 and n11272 n11283_not ; n11285
g11030 and n11284_not n11285_not ; n11286
g11031 and n10918_not n11286 ; n11287
g11032 and n10918 n11286_not ; n11288
g11033 and n11287_not n11288_not ; n11289
g11034 and n11121_not n11289 ; n11290
g11035 and n11121 n11289_not ; n11291
g11036 and n11290_not n11291_not ; n11292
g11037 and n11110_not n11292 ; n11293
g11038 and n11110 n11292_not ; n11294
g11039 and n11293_not n11294_not ; n11295
g11040 and b[33] n2539 ; n11296
g11041 and b[31] n2685 ; n11297
g11042 and b[32] n2534 ; n11298
g11043 and n11297_not n11298_not ; n11299
g11044 and n11296_not n11299 ; n11300
g11045 and n2542 n4223 ; n11301
g11046 and n11300 n11301_not ; n11302
g11047 and a[26] n11302_not ; n11303
g11048 and a[26] n11303_not ; n11304
g11049 and n11302_not n11303_not ; n11305
g11050 and n11304_not n11305_not ; n11306
g11051 and n11295 n11306_not ; n11307
g11052 and n11295 n11307_not ; n11308
g11053 and n11306_not n11307_not ; n11309
g11054 and n11308_not n11309_not ; n11310
g11055 and n11109_not n11310 ; n11311
g11056 and n11109 n11310_not ; n11312
g11057 and n11311_not n11312_not ; n11313
g11058 and b[36] n2048 ; n11314
g11059 and b[34] n2198 ; n11315
g11060 and b[35] n2043 ; n11316
g11061 and n11315_not n11316_not ; n11317
g11062 and n11314_not n11317 ; n11318
g11063 and n2051 n4922 ; n11319
g11064 and n11318 n11319_not ; n11320
g11065 and a[23] n11320_not ; n11321
g11066 and a[23] n11321_not ; n11322
g11067 and n11320_not n11321_not ; n11323
g11068 and n11322_not n11323_not ; n11324
g11069 and n11313_not n11324_not ; n11325
g11070 and n11313 n11324 ; n11326
g11071 and n11325_not n11326_not ; n11327
g11072 and n11108 n11327_not ; n11328
g11073 and n11108_not n11327 ; n11329
g11074 and n11328_not n11329_not ; n11330
g11075 and b[39] n1627 ; n11331
g11076 and b[37] n1763 ; n11332
g11077 and b[38] n1622 ; n11333
g11078 and n11332_not n11333_not ; n11334
g11079 and n11331_not n11334 ; n11335
g11080 and n1630 n5451 ; n11336
g11081 and n11335 n11336_not ; n11337
g11082 and a[20] n11337_not ; n11338
g11083 and a[20] n11338_not ; n11339
g11084 and n11337_not n11338_not ; n11340
g11085 and n11339_not n11340_not ; n11341
g11086 and n11330 n11341_not ; n11342
g11087 and n11330 n11342_not ; n11343
g11088 and n11341_not n11342_not ; n11344
g11089 and n11343_not n11344_not ; n11345
g11090 and n10963_not n10969_not ; n11346
g11091 and n11345 n11346 ; n11347
g11092 and n11345_not n11346_not ; n11348
g11093 and n11347_not n11348_not ; n11349
g11094 and b[42] n1302 ; n11350
g11095 and b[40] n1391 ; n11351
g11096 and b[41] n1297 ; n11352
g11097 and n11351_not n11352_not ; n11353
g11098 and n11350_not n11353 ; n11354
g11099 and n1305 n6489 ; n11355
g11100 and n11354 n11355_not ; n11356
g11101 and a[17] n11356_not ; n11357
g11102 and a[17] n11357_not ; n11358
g11103 and n11356_not n11357_not ; n11359
g11104 and n11358_not n11359_not ; n11360
g11105 and n11349_not n11360 ; n11361
g11106 and n11349 n11360_not ; n11362
g11107 and n11361_not n11362_not ; n11363
g11108 and n11107_not n11363 ; n11364
g11109 and n11107 n11363_not ; n11365
g11110 and n11364_not n11365_not ; n11366
g11111 and n11106_not n11366 ; n11367
g11112 and n11106_not n11367_not ; n11368
g11113 and n11366 n11367_not ; n11369
g11114 and n11368_not n11369_not ; n11370
g11115 and n11006_not n11370_not ; n11371
g11116 and n11006 n11369_not ; n11372
g11117 and n11368_not n11372 ; n11373
g11118 and n11371_not n11373_not ; n11374
g11119 and n11095_not n11374 ; n11375
g11120 and n11095_not n11375_not ; n11376
g11121 and n11374 n11375_not ; n11377
g11122 and n11376_not n11377_not ; n11378
g11123 and n11084_not n11378_not ; n11379
g11124 and n11084 n11377_not ; n11380
g11125 and n11376_not n11380 ; n11381
g11126 and n11379_not n11381_not ; n11382
g11127 and n11083_not n11382 ; n11383
g11128 and n11083_not n11383_not ; n11384
g11129 and n11382 n11383_not ; n11385
g11130 and n11384_not n11385_not ; n11386
g11131 and n11072_not n11386_not ; n11387
g11132 and n11072 n11385_not ; n11388
g11133 and n11384_not n11388 ; n11389
g11134 and n11387_not n11389_not ; n11390
g11135 and n11071_not n11390 ; n11391
g11136 and n11071_not n11391_not ; n11392
g11137 and n11390 n11391_not ; n11393
g11138 and n11392_not n11393_not ; n11394
g11139 and n11060_not n11394_not ; n11395
g11140 and n11060_not n11395_not ; n11396
g11141 and n11394_not n11395_not ; n11397
g11142 and n11396_not n11397_not ; n11398
g11143 and b[57] n266 ; n11399
g11144 and b[55] n284 ; n11400
g11145 and b[56] n261 ; n11401
g11146 and n11400_not n11401_not ; n11402
g11147 and n11399_not n11402 ; n11403
g11148 and n10704_not n10706_not ; n11404
g11149 and b[56]_not b[57]_not ; n11405
g11150 and b[56] b[57] ; n11406
g11151 and n11405_not n11406_not ; n11407
g11152 and n11404_not n11407 ; n11408
g11153 and n11404 n11407_not ; n11409
g11154 and n11408_not n11409_not ; n11410
g11155 and n269 n11410 ; n11411
g11156 and n11403 n11411_not ; n11412
g11157 and a[2] n11412_not ; n11413
g11158 and a[2] n11413_not ; n11414
g11159 and n11412_not n11413_not ; n11415
g11160 and n11414_not n11415_not ; n11416
g11161 and n11398_not n11416_not ; n11417
g11162 and n11398_not n11417_not ; n11418
g11163 and n11416_not n11417_not ; n11419
g11164 and n11418_not n11419_not ; n11420
g11165 and n11052_not n11057_not ; n11421
g11166 and n11420_not n11421_not ; n11422
g11167 and n11420 n11421 ; n11423
g11168 and n11422_not n11423_not ; f[57]
g11169 and b[58] n266 ; n11425
g11170 and b[56] n284 ; n11426
g11171 and b[57] n261 ; n11427
g11172 and n11426_not n11427_not ; n11428
g11173 and n11425_not n11428 ; n11429
g11174 and n11406_not n11408_not ; n11430
g11175 and b[57]_not b[58]_not ; n11431
g11176 and b[57] b[58] ; n11432
g11177 and n11431_not n11432_not ; n11433
g11178 and n11430_not n11433 ; n11434
g11179 and n11430 n11433_not ; n11435
g11180 and n11434_not n11435_not ; n11436
g11181 and n269 n11436 ; n11437
g11182 and n11429 n11437_not ; n11438
g11183 and a[2] n11438_not ; n11439
g11184 and a[2] n11439_not ; n11440
g11185 and n11438_not n11439_not ; n11441
g11186 and n11440_not n11441_not ; n11442
g11187 and n11391_not n11395_not ; n11443
g11188 and b[55] n362 ; n11444
g11189 and b[53] n403 ; n11445
g11190 and b[54] n357 ; n11446
g11191 and n11445_not n11446_not ; n11447
g11192 and n11444_not n11447 ; n11448
g11193 and n365 n10684 ; n11449
g11194 and n11448 n11449_not ; n11450
g11195 and a[5] n11450_not ; n11451
g11196 and a[5] n11451_not ; n11452
g11197 and n11450_not n11451_not ; n11453
g11198 and n11452_not n11453_not ; n11454
g11199 and n11383_not n11387_not ; n11455
g11200 and b[52] n511 ; n11456
g11201 and b[50] n541 ; n11457
g11202 and b[51] n506 ; n11458
g11203 and n11457_not n11458_not ; n11459
g11204 and n11456_not n11459 ; n11460
g11205 and n514 n9628 ; n11461
g11206 and n11460 n11461_not ; n11462
g11207 and a[8] n11462_not ; n11463
g11208 and a[8] n11463_not ; n11464
g11209 and n11462_not n11463_not ; n11465
g11210 and n11464_not n11465_not ; n11466
g11211 and n11375_not n11379_not ; n11467
g11212 and b[49] n700 ; n11468
g11213 and b[47] n767 ; n11469
g11214 and b[48] n695 ; n11470
g11215 and n11469_not n11470_not ; n11471
g11216 and n11468_not n11471 ; n11472
g11217 and n703 n8625 ; n11473
g11218 and n11472 n11473_not ; n11474
g11219 and a[11] n11474_not ; n11475
g11220 and a[11] n11475_not ; n11476
g11221 and n11474_not n11475_not ; n11477
g11222 and n11476_not n11477_not ; n11478
g11223 and n11367_not n11371_not ; n11479
g11224 and n11362_not n11364_not ; n11480
g11225 and n11290_not n11293_not ; n11481
g11226 and n11285_not n11287_not ; n11482
g11227 and n11240_not n11244_not ; n11483
g11228 and n11229_not n11231_not ; n11484
g11229 and b[10] n8362 ; n11485
g11230 and b[8] n8715 ; n11486
g11231 and b[9] n8357 ; n11487
g11232 and n11486_not n11487_not ; n11488
g11233 and n11485_not n11488 ; n11489
g11234 and n738 n8365 ; n11490
g11235 and n11489 n11490_not ; n11491
g11236 and a[50] n11491_not ; n11492
g11237 and a[50] n11492_not ; n11493
g11238 and n11491_not n11492_not ; n11494
g11239 and n11493_not n11494_not ; n11495
g11240 and n10826_not n11207_not ; n11496
g11241 and n11204_not n11496_not ; n11497
g11242 and b[7] n9339 ; n11498
g11243 and b[5] n9732 ; n11499
g11244 and b[6] n9334 ; n11500
g11245 and n11499_not n11500_not ; n11501
g11246 and n11498_not n11501 ; n11502
g11247 and n484 n9342 ; n11503
g11248 and n11502 n11503_not ; n11504
g11249 and a[53] n11504_not ; n11505
g11250 and a[53] n11505_not ; n11506
g11251 and n11504_not n11505_not ; n11507
g11252 and n11506_not n11507_not ; n11508
g11253 and n10808 n11186 ; n11509
g11254 and n11201_not n11509_not ; n11510
g11255 and b[4] n10426 ; n11511
g11256 and b[2] n10796 ; n11512
g11257 and b[3] n10421 ; n11513
g11258 and n11512_not n11513_not ; n11514
g11259 and n11511_not n11514 ; n11515
g11260 and n346 n10429 ; n11516
g11261 and n11515 n11516_not ; n11517
g11262 and a[56] n11517_not ; n11518
g11263 and a[56] n11518_not ; n11519
g11264 and n11517_not n11518_not ; n11520
g11265 and n11519_not n11520_not ; n11521
g11266 and a[59] n11186_not ; n11522
g11267 and a[57]_not a[58] ; n11523
g11268 and a[57] a[58]_not ; n11524
g11269 and n11523_not n11524_not ; n11525
g11270 and n11185 n11525_not ; n11526
g11271 and b[0] n11526 ; n11527
g11272 and a[58]_not a[59] ; n11528
g11273 and a[58] a[59]_not ; n11529
g11274 and n11528_not n11529_not ; n11530
g11275 and n11185_not n11530 ; n11531
g11276 and b[1] n11531 ; n11532
g11277 and n11527_not n11532_not ; n11533
g11278 and n11185_not n11530_not ; n11534
g11279 and n272_not n11534 ; n11535
g11280 and n11533 n11535_not ; n11536
g11281 and a[59] n11536_not ; n11537
g11282 and a[59] n11537_not ; n11538
g11283 and n11536_not n11537_not ; n11539
g11284 and n11538_not n11539_not ; n11540
g11285 and n11522 n11540_not ; n11541
g11286 and n11522_not n11540 ; n11542
g11287 and n11541_not n11542_not ; n11543
g11288 and n11521 n11543_not ; n11544
g11289 and n11521_not n11543 ; n11545
g11290 and n11544_not n11545_not ; n11546
g11291 and n11510_not n11546 ; n11547
g11292 and n11510 n11546_not ; n11548
g11293 and n11547_not n11548_not ; n11549
g11294 and n11508 n11549_not ; n11550
g11295 and n11508_not n11549 ; n11551
g11296 and n11550_not n11551_not ; n11552
g11297 and n11497_not n11552 ; n11553
g11298 and n11497 n11552_not ; n11554
g11299 and n11553_not n11554_not ; n11555
g11300 and n11495_not n11555 ; n11556
g11301 and n11555 n11556_not ; n11557
g11302 and n11495_not n11556_not ; n11558
g11303 and n11557_not n11558_not ; n11559
g11304 and n11222_not n11225_not ; n11560
g11305 and n11559 n11560 ; n11561
g11306 and n11559_not n11560_not ; n11562
g11307 and n11561_not n11562_not ; n11563
g11308 and b[13] n7446 ; n11564
g11309 and b[11] n7787 ; n11565
g11310 and b[12] n7441 ; n11566
g11311 and n11565_not n11566_not ; n11567
g11312 and n11564_not n11567 ; n11568
g11313 and n1008 n7449 ; n11569
g11314 and n11568 n11569_not ; n11570
g11315 and a[47] n11570_not ; n11571
g11316 and a[47] n11571_not ; n11572
g11317 and n11570_not n11571_not ; n11573
g11318 and n11572_not n11573_not ; n11574
g11319 and n11563 n11574_not ; n11575
g11320 and n11563_not n11574 ; n11576
g11321 and n11484_not n11576_not ; n11577
g11322 and n11575_not n11577 ; n11578
g11323 and n11484_not n11578_not ; n11579
g11324 and n11575_not n11578_not ; n11580
g11325 and n11576_not n11580 ; n11581
g11326 and n11579_not n11581_not ; n11582
g11327 and b[16] n6595 ; n11583
g11328 and b[14] n6902 ; n11584
g11329 and b[15] n6590 ; n11585
g11330 and n11584_not n11585_not ; n11586
g11331 and n11583_not n11586 ; n11587
g11332 and n1237 n6598 ; n11588
g11333 and n11587 n11588_not ; n11589
g11334 and a[44] n11589_not ; n11590
g11335 and a[44] n11590_not ; n11591
g11336 and n11589_not n11590_not ; n11592
g11337 and n11591_not n11592_not ; n11593
g11338 and n11582_not n11593_not ; n11594
g11339 and n11582_not n11594_not ; n11595
g11340 and n11593_not n11594_not ; n11596
g11341 and n11595_not n11596_not ; n11597
g11342 and n11234_not n11237_not ; n11598
g11343 and n11597 n11598 ; n11599
g11344 and n11597_not n11598_not ; n11600
g11345 and n11599_not n11600_not ; n11601
g11346 and b[19] n5777 ; n11602
g11347 and b[17] n6059 ; n11603
g11348 and b[18] n5772 ; n11604
g11349 and n11603_not n11604_not ; n11605
g11350 and n11602_not n11605 ; n11606
g11351 and n1708 n5780 ; n11607
g11352 and n11606 n11607_not ; n11608
g11353 and a[41] n11608_not ; n11609
g11354 and a[41] n11609_not ; n11610
g11355 and n11608_not n11609_not ; n11611
g11356 and n11610_not n11611_not ; n11612
g11357 and n11601 n11612_not ; n11613
g11358 and n11601_not n11612 ; n11614
g11359 and n11483_not n11614_not ; n11615
g11360 and n11613_not n11615 ; n11616
g11361 and n11483_not n11616_not ; n11617
g11362 and n11613_not n11616_not ; n11618
g11363 and n11614_not n11618 ; n11619
g11364 and n11617_not n11619_not ; n11620
g11365 and b[22] n5035 ; n11621
g11366 and b[20] n5277 ; n11622
g11367 and b[21] n5030 ; n11623
g11368 and n11622_not n11623_not ; n11624
g11369 and n11621_not n11624 ; n11625
g11370 and n2145 n5038 ; n11626
g11371 and n11625 n11626_not ; n11627
g11372 and a[38] n11627_not ; n11628
g11373 and a[38] n11628_not ; n11629
g11374 and n11627_not n11628_not ; n11630
g11375 and n11629_not n11630_not ; n11631
g11376 and n11620_not n11631_not ; n11632
g11377 and n11620_not n11632_not ; n11633
g11378 and n11631_not n11632_not ; n11634
g11379 and n11633_not n11634_not ; n11635
g11380 and n11248_not n11251_not ; n11636
g11381 and n11635 n11636 ; n11637
g11382 and n11635_not n11636_not ; n11638
g11383 and n11637_not n11638_not ; n11639
g11384 and b[25] n4287 ; n11640
g11385 and b[23] n4532 ; n11641
g11386 and b[24] n4282 ; n11642
g11387 and n11641_not n11642_not ; n11643
g11388 and n11640_not n11643 ; n11644
g11389 and n2485 n4290 ; n11645
g11390 and n11644 n11645_not ; n11646
g11391 and a[35] n11646_not ; n11647
g11392 and a[35] n11647_not ; n11648
g11393 and n11646_not n11647_not ; n11649
g11394 and n11648_not n11649_not ; n11650
g11395 and n11639 n11650_not ; n11651
g11396 and n11639 n11651_not ; n11652
g11397 and n11650_not n11651_not ; n11653
g11398 and n11652_not n11653_not ; n11654
g11399 and n11265_not n11271_not ; n11655
g11400 and n11654 n11655 ; n11656
g11401 and n11654_not n11655_not ; n11657
g11402 and n11656_not n11657_not ; n11658
g11403 and b[28] n3638 ; n11659
g11404 and b[26] n3843 ; n11660
g11405 and b[27] n3633 ; n11661
g11406 and n11660_not n11661_not ; n11662
g11407 and n11659_not n11662 ; n11663
g11408 and n3189 n3641 ; n11664
g11409 and n11663 n11664_not ; n11665
g11410 and a[32] n11665_not ; n11666
g11411 and a[32] n11666_not ; n11667
g11412 and n11665_not n11666_not ; n11668
g11413 and n11667_not n11668_not ; n11669
g11414 and n11658 n11669_not ; n11670
g11415 and n11658 n11670_not ; n11671
g11416 and n11669_not n11670_not ; n11672
g11417 and n11671_not n11672_not ; n11673
g11418 and n11482_not n11673 ; n11674
g11419 and n11482 n11673_not ; n11675
g11420 and n11674_not n11675_not ; n11676
g11421 and b[31] n3050 ; n11677
g11422 and b[29] n3243 ; n11678
g11423 and b[30] n3045 ; n11679
g11424 and n11678_not n11679_not ; n11680
g11425 and n11677_not n11680 ; n11681
g11426 and n3053 n3796 ; n11682
g11427 and n11681 n11682_not ; n11683
g11428 and a[29] n11683_not ; n11684
g11429 and a[29] n11684_not ; n11685
g11430 and n11683_not n11684_not ; n11686
g11431 and n11685_not n11686_not ; n11687
g11432 and n11676_not n11687_not ; n11688
g11433 and n11676 n11687 ; n11689
g11434 and n11688_not n11689_not ; n11690
g11435 and n11481 n11690_not ; n11691
g11436 and n11481_not n11690 ; n11692
g11437 and n11691_not n11692_not ; n11693
g11438 and b[34] n2539 ; n11694
g11439 and b[32] n2685 ; n11695
g11440 and b[33] n2534 ; n11696
g11441 and n11695_not n11696_not ; n11697
g11442 and n11694_not n11697 ; n11698
g11443 and n2542 n4466 ; n11699
g11444 and n11698 n11699_not ; n11700
g11445 and a[26] n11700_not ; n11701
g11446 and a[26] n11701_not ; n11702
g11447 and n11700_not n11701_not ; n11703
g11448 and n11702_not n11703_not ; n11704
g11449 and n11693 n11704_not ; n11705
g11450 and n11693 n11705_not ; n11706
g11451 and n11704_not n11705_not ; n11707
g11452 and n11706_not n11707_not ; n11708
g11453 and n11109_not n11310_not ; n11709
g11454 and n11307_not n11709_not ; n11710
g11455 and n11708 n11710 ; n11711
g11456 and n11708_not n11710_not ; n11712
g11457 and n11711_not n11712_not ; n11713
g11458 and b[37] n2048 ; n11714
g11459 and b[35] n2198 ; n11715
g11460 and b[36] n2043 ; n11716
g11461 and n11715_not n11716_not ; n11717
g11462 and n11714_not n11717 ; n11718
g11463 and n2051 n5181 ; n11719
g11464 and n11718 n11719_not ; n11720
g11465 and a[23] n11720_not ; n11721
g11466 and a[23] n11721_not ; n11722
g11467 and n11720_not n11721_not ; n11723
g11468 and n11722_not n11723_not ; n11724
g11469 and n11713 n11724_not ; n11725
g11470 and n11713 n11725_not ; n11726
g11471 and n11724_not n11725_not ; n11727
g11472 and n11726_not n11727_not ; n11728
g11473 and n11325_not n11329_not ; n11729
g11474 and n11728 n11729 ; n11730
g11475 and n11728_not n11729_not ; n11731
g11476 and n11730_not n11731_not ; n11732
g11477 and b[40] n1627 ; n11733
g11478 and b[38] n1763 ; n11734
g11479 and b[39] n1622 ; n11735
g11480 and n11734_not n11735_not ; n11736
g11481 and n11733_not n11736 ; n11737
g11482 and n1630 n5955 ; n11738
g11483 and n11737 n11738_not ; n11739
g11484 and a[20] n11739_not ; n11740
g11485 and a[20] n11740_not ; n11741
g11486 and n11739_not n11740_not ; n11742
g11487 and n11741_not n11742_not ; n11743
g11488 and n11732 n11743_not ; n11744
g11489 and n11732 n11744_not ; n11745
g11490 and n11743_not n11744_not ; n11746
g11491 and n11745_not n11746_not ; n11747
g11492 and n11342_not n11348_not ; n11748
g11493 and n11747 n11748 ; n11749
g11494 and n11747_not n11748_not ; n11750
g11495 and n11749_not n11750_not ; n11751
g11496 and b[43] n1302 ; n11752
g11497 and b[41] n1391 ; n11753
g11498 and b[42] n1297 ; n11754
g11499 and n11753_not n11754_not ; n11755
g11500 and n11752_not n11755 ; n11756
g11501 and n1305 n6515 ; n11757
g11502 and n11756 n11757_not ; n11758
g11503 and a[17] n11758_not ; n11759
g11504 and a[17] n11759_not ; n11760
g11505 and n11758_not n11759_not ; n11761
g11506 and n11760_not n11761_not ; n11762
g11507 and n11751 n11762_not ; n11763
g11508 and n11751_not n11762 ; n11764
g11509 and n11480_not n11764_not ; n11765
g11510 and n11763_not n11765 ; n11766
g11511 and n11480_not n11766_not ; n11767
g11512 and n11763_not n11766_not ; n11768
g11513 and n11764_not n11768 ; n11769
g11514 and n11767_not n11769_not ; n11770
g11515 and b[46] n951 ; n11771
g11516 and b[44] n1056 ; n11772
g11517 and b[45] n946 ; n11773
g11518 and n11772_not n11773_not ; n11774
g11519 and n11771_not n11774 ; n11775
g11520 and n954 n7677 ; n11776
g11521 and n11775 n11776_not ; n11777
g11522 and a[14] n11777_not ; n11778
g11523 and a[14] n11778_not ; n11779
g11524 and n11777_not n11778_not ; n11780
g11525 and n11779_not n11780_not ; n11781
g11526 and n11770 n11781 ; n11782
g11527 and n11770_not n11781_not ; n11783
g11528 and n11782_not n11783_not ; n11784
g11529 and n11479_not n11784 ; n11785
g11530 and n11479 n11784_not ; n11786
g11531 and n11785_not n11786_not ; n11787
g11532 and n11478 n11787_not ; n11788
g11533 and n11478_not n11787 ; n11789
g11534 and n11788_not n11789_not ; n11790
g11535 and n11467_not n11790 ; n11791
g11536 and n11467 n11790_not ; n11792
g11537 and n11791_not n11792_not ; n11793
g11538 and n11466 n11793_not ; n11794
g11539 and n11466_not n11793 ; n11795
g11540 and n11794_not n11795_not ; n11796
g11541 and n11455_not n11796 ; n11797
g11542 and n11455 n11796_not ; n11798
g11543 and n11797_not n11798_not ; n11799
g11544 and n11454 n11799_not ; n11800
g11545 and n11454_not n11799 ; n11801
g11546 and n11800_not n11801_not ; n11802
g11547 and n11443_not n11802 ; n11803
g11548 and n11443 n11802_not ; n11804
g11549 and n11803_not n11804_not ; n11805
g11550 and n11442_not n11805 ; n11806
g11551 and n11805 n11806_not ; n11807
g11552 and n11442_not n11806_not ; n11808
g11553 and n11807_not n11808_not ; n11809
g11554 and n11417_not n11422_not ; n11810
g11555 and n11809_not n11810_not ; n11811
g11556 and n11809 n11810 ; n11812
g11557 and n11811_not n11812_not ; f[58]
g11558 and n11806_not n11811_not ; n11814
g11559 and n11801_not n11803_not ; n11815
g11560 and n11795_not n11797_not ; n11816
g11561 and b[53] n511 ; n11817
g11562 and b[51] n541 ; n11818
g11563 and b[52] n506 ; n11819
g11564 and n11818_not n11819_not ; n11820
g11565 and n11817_not n11820 ; n11821
g11566 and n514 n9972 ; n11822
g11567 and n11821 n11822_not ; n11823
g11568 and a[8] n11823_not ; n11824
g11569 and a[8] n11824_not ; n11825
g11570 and n11823_not n11824_not ; n11826
g11571 and n11825_not n11826_not ; n11827
g11572 and n11789_not n11791_not ; n11828
g11573 and b[50] n700 ; n11829
g11574 and b[48] n767 ; n11830
g11575 and b[49] n695 ; n11831
g11576 and n11830_not n11831_not ; n11832
g11577 and n11829_not n11832 ; n11833
g11578 and n703 n8949 ; n11834
g11579 and n11833 n11834_not ; n11835
g11580 and a[11] n11835_not ; n11836
g11581 and a[11] n11836_not ; n11837
g11582 and n11835_not n11836_not ; n11838
g11583 and n11837_not n11838_not ; n11839
g11584 and n11783_not n11785_not ; n11840
g11585 and n11744_not n11750_not ; n11841
g11586 and b[35] n2539 ; n11842
g11587 and b[33] n2685 ; n11843
g11588 and b[34] n2534 ; n11844
g11589 and n11843_not n11844_not ; n11845
g11590 and n11842_not n11845 ; n11846
g11591 and n2542 n4696 ; n11847
g11592 and n11846 n11847_not ; n11848
g11593 and a[26] n11848_not ; n11849
g11594 and a[26] n11849_not ; n11850
g11595 and n11848_not n11849_not ; n11851
g11596 and n11850_not n11851_not ; n11852
g11597 and n11688_not n11692_not ; n11853
g11598 and n11482_not n11673_not ; n11854
g11599 and n11670_not n11854_not ; n11855
g11600 and n11632_not n11638_not ; n11856
g11601 and n11594_not n11600_not ; n11857
g11602 and b[17] n6595 ; n11858
g11603 and b[15] n6902 ; n11859
g11604 and b[16] n6590 ; n11860
g11605 and n11859_not n11860_not ; n11861
g11606 and n11858_not n11861 ; n11862
g11607 and n1356 n6598 ; n11863
g11608 and n11862 n11863_not ; n11864
g11609 and a[44] n11864_not ; n11865
g11610 and a[44] n11865_not ; n11866
g11611 and n11864_not n11865_not ; n11867
g11612 and n11866_not n11867_not ; n11868
g11613 and b[14] n7446 ; n11869
g11614 and b[12] n7787 ; n11870
g11615 and b[13] n7441 ; n11871
g11616 and n11870_not n11871_not ; n11872
g11617 and n11869_not n11872 ; n11873
g11618 and n1034 n7449 ; n11874
g11619 and n11873 n11874_not ; n11875
g11620 and a[47] n11875_not ; n11876
g11621 and a[47] n11876_not ; n11877
g11622 and n11875_not n11876_not ; n11878
g11623 and n11877_not n11878_not ; n11879
g11624 and n11556_not n11562_not ; n11880
g11625 and b[11] n8362 ; n11881
g11626 and b[9] n8715 ; n11882
g11627 and b[10] n8357 ; n11883
g11628 and n11882_not n11883_not ; n11884
g11629 and n11881_not n11884 ; n11885
g11630 and n818 n8365 ; n11886
g11631 and n11885 n11886_not ; n11887
g11632 and a[50] n11887_not ; n11888
g11633 and a[50] n11888_not ; n11889
g11634 and n11887_not n11888_not ; n11890
g11635 and n11889_not n11890_not ; n11891
g11636 and n11551_not n11553_not ; n11892
g11637 and n11545_not n11547_not ; n11893
g11638 and b[2] n11531 ; n11894
g11639 and n11185 n11530_not ; n11895
g11640 and n11525 n11895 ; n11896
g11641 and b[0] n11896 ; n11897
g11642 and b[1] n11526 ; n11898
g11643 and n11897_not n11898_not ; n11899
g11644 and n11894_not n11899 ; n11900
g11645 and n296 n11534 ; n11901
g11646 and n11900 n11901_not ; n11902
g11647 and a[59] n11902_not ; n11903
g11648 and a[59] n11903_not ; n11904
g11649 and n11902_not n11903_not ; n11905
g11650 and n11904_not n11905_not ; n11906
g11651 and n11541_not n11906 ; n11907
g11652 and n11541 n11906_not ; n11908
g11653 and n11907_not n11908_not ; n11909
g11654 and b[5] n10426 ; n11910
g11655 and b[3] n10796 ; n11911
g11656 and b[4] n10421 ; n11912
g11657 and n11911_not n11912_not ; n11913
g11658 and n11910_not n11913 ; n11914
g11659 and n394 n10429 ; n11915
g11660 and n11914 n11915_not ; n11916
g11661 and a[56] n11916_not ; n11917
g11662 and a[56] n11917_not ; n11918
g11663 and n11916_not n11917_not ; n11919
g11664 and n11918_not n11919_not ; n11920
g11665 and n11909 n11920_not ; n11921
g11666 and n11909_not n11920 ; n11922
g11667 and n11893_not n11922_not ; n11923
g11668 and n11921_not n11923 ; n11924
g11669 and n11893_not n11924_not ; n11925
g11670 and n11921_not n11924_not ; n11926
g11671 and n11922_not n11926 ; n11927
g11672 and n11925_not n11927_not ; n11928
g11673 and b[8] n9339 ; n11929
g11674 and b[6] n9732 ; n11930
g11675 and b[7] n9334 ; n11931
g11676 and n11930_not n11931_not ; n11932
g11677 and n11929_not n11932 ; n11933
g11678 and n585 n9342 ; n11934
g11679 and n11933 n11934_not ; n11935
g11680 and a[53] n11935_not ; n11936
g11681 and a[53] n11936_not ; n11937
g11682 and n11935_not n11936_not ; n11938
g11683 and n11937_not n11938_not ; n11939
g11684 and n11928 n11939 ; n11940
g11685 and n11928_not n11939_not ; n11941
g11686 and n11940_not n11941_not ; n11942
g11687 and n11892_not n11942 ; n11943
g11688 and n11892 n11942_not ; n11944
g11689 and n11943_not n11944_not ; n11945
g11690 and n11891 n11945_not ; n11946
g11691 and n11891_not n11945 ; n11947
g11692 and n11946_not n11947_not ; n11948
g11693 and n11880_not n11948 ; n11949
g11694 and n11880 n11948_not ; n11950
g11695 and n11949_not n11950_not ; n11951
g11696 and n11879_not n11951 ; n11952
g11697 and n11951 n11952_not ; n11953
g11698 and n11879_not n11952_not ; n11954
g11699 and n11953_not n11954_not ; n11955
g11700 and n11580_not n11955_not ; n11956
g11701 and n11580 n11955 ; n11957
g11702 and n11956_not n11957_not ; n11958
g11703 and n11868_not n11958 ; n11959
g11704 and n11868_not n11959_not ; n11960
g11705 and n11958 n11959_not ; n11961
g11706 and n11960_not n11961_not ; n11962
g11707 and n11857_not n11962_not ; n11963
g11708 and n11857_not n11963_not ; n11964
g11709 and n11962_not n11963_not ; n11965
g11710 and n11964_not n11965_not ; n11966
g11711 and b[20] n5777 ; n11967
g11712 and b[18] n6059 ; n11968
g11713 and b[19] n5772 ; n11969
g11714 and n11968_not n11969_not ; n11970
g11715 and n11967_not n11970 ; n11971
g11716 and n1846 n5780 ; n11972
g11717 and n11971 n11972_not ; n11973
g11718 and a[41] n11973_not ; n11974
g11719 and a[41] n11974_not ; n11975
g11720 and n11973_not n11974_not ; n11976
g11721 and n11975_not n11976_not ; n11977
g11722 and n11966_not n11977_not ; n11978
g11723 and n11966_not n11978_not ; n11979
g11724 and n11977_not n11978_not ; n11980
g11725 and n11979_not n11980_not ; n11981
g11726 and n11618_not n11981 ; n11982
g11727 and n11618 n11981_not ; n11983
g11728 and n11982_not n11983_not ; n11984
g11729 and b[23] n5035 ; n11985
g11730 and b[21] n5277 ; n11986
g11731 and b[22] n5030 ; n11987
g11732 and n11986_not n11987_not ; n11988
g11733 and n11985_not n11988 ; n11989
g11734 and n2300 n5038 ; n11990
g11735 and n11989 n11990_not ; n11991
g11736 and a[38] n11991_not ; n11992
g11737 and a[38] n11992_not ; n11993
g11738 and n11991_not n11992_not ; n11994
g11739 and n11993_not n11994_not ; n11995
g11740 and n11984_not n11995_not ; n11996
g11741 and n11984 n11995 ; n11997
g11742 and n11996_not n11997_not ; n11998
g11743 and n11856 n11998_not ; n11999
g11744 and n11856_not n11998 ; n12000
g11745 and n11999_not n12000_not ; n12001
g11746 and b[26] n4287 ; n12002
g11747 and b[24] n4532 ; n12003
g11748 and b[25] n4282 ; n12004
g11749 and n12003_not n12004_not ; n12005
g11750 and n12002_not n12005 ; n12006
g11751 and n2813 n4290 ; n12007
g11752 and n12006 n12007_not ; n12008
g11753 and a[35] n12008_not ; n12009
g11754 and a[35] n12009_not ; n12010
g11755 and n12008_not n12009_not ; n12011
g11756 and n12010_not n12011_not ; n12012
g11757 and n12001 n12012_not ; n12013
g11758 and n12001 n12013_not ; n12014
g11759 and n12012_not n12013_not ; n12015
g11760 and n12014_not n12015_not ; n12016
g11761 and n11651_not n11657_not ; n12017
g11762 and n12016 n12017 ; n12018
g11763 and n12016_not n12017_not ; n12019
g11764 and n12018_not n12019_not ; n12020
g11765 and b[29] n3638 ; n12021
g11766 and b[27] n3843 ; n12022
g11767 and b[28] n3633 ; n12023
g11768 and n12022_not n12023_not ; n12024
g11769 and n12021_not n12024 ; n12025
g11770 and n3383 n3641 ; n12026
g11771 and n12025 n12026_not ; n12027
g11772 and a[32] n12027_not ; n12028
g11773 and a[32] n12028_not ; n12029
g11774 and n12027_not n12028_not ; n12030
g11775 and n12029_not n12030_not ; n12031
g11776 and n12020 n12031_not ; n12032
g11777 and n12020_not n12031 ; n12033
g11778 and n11855_not n12033_not ; n12034
g11779 and n12032_not n12034 ; n12035
g11780 and n11855_not n12035_not ; n12036
g11781 and n12032_not n12035_not ; n12037
g11782 and n12033_not n12037 ; n12038
g11783 and n12036_not n12038_not ; n12039
g11784 and b[32] n3050 ; n12040
g11785 and b[30] n3243 ; n12041
g11786 and b[31] n3045 ; n12042
g11787 and n12041_not n12042_not ; n12043
g11788 and n12040_not n12043 ; n12044
g11789 and n3053 n4013 ; n12045
g11790 and n12044 n12045_not ; n12046
g11791 and a[29] n12046_not ; n12047
g11792 and a[29] n12047_not ; n12048
g11793 and n12046_not n12047_not ; n12049
g11794 and n12048_not n12049_not ; n12050
g11795 and n12039 n12050 ; n12051
g11796 and n12039_not n12050_not ; n12052
g11797 and n12051_not n12052_not ; n12053
g11798 and n11853_not n12053 ; n12054
g11799 and n11853 n12053_not ; n12055
g11800 and n12054_not n12055_not ; n12056
g11801 and n11852_not n12056 ; n12057
g11802 and n12056 n12057_not ; n12058
g11803 and n11852_not n12057_not ; n12059
g11804 and n12058_not n12059_not ; n12060
g11805 and n11705_not n11712_not ; n12061
g11806 and n12060 n12061 ; n12062
g11807 and n12060_not n12061_not ; n12063
g11808 and n12062_not n12063_not ; n12064
g11809 and b[38] n2048 ; n12065
g11810 and b[36] n2198 ; n12066
g11811 and b[37] n2043 ; n12067
g11812 and n12066_not n12067_not ; n12068
g11813 and n12065_not n12068 ; n12069
g11814 and n2051 n5205 ; n12070
g11815 and n12069 n12070_not ; n12071
g11816 and a[23] n12071_not ; n12072
g11817 and a[23] n12072_not ; n12073
g11818 and n12071_not n12072_not ; n12074
g11819 and n12073_not n12074_not ; n12075
g11820 and n12064 n12075_not ; n12076
g11821 and n12064 n12076_not ; n12077
g11822 and n12075_not n12076_not ; n12078
g11823 and n12077_not n12078_not ; n12079
g11824 and n11725_not n11731_not ; n12080
g11825 and n12079 n12080 ; n12081
g11826 and n12079_not n12080_not ; n12082
g11827 and n12081_not n12082_not ; n12083
g11828 and b[41] n1627 ; n12084
g11829 and b[39] n1763 ; n12085
g11830 and b[40] n1622 ; n12086
g11831 and n12085_not n12086_not ; n12087
g11832 and n12084_not n12087 ; n12088
g11833 and n1630 n6219 ; n12089
g11834 and n12088 n12089_not ; n12090
g11835 and a[20] n12090_not ; n12091
g11836 and a[20] n12091_not ; n12092
g11837 and n12090_not n12091_not ; n12093
g11838 and n12092_not n12093_not ; n12094
g11839 and n12083 n12094_not ; n12095
g11840 and n12083_not n12094 ; n12096
g11841 and n11841_not n12096_not ; n12097
g11842 and n12095_not n12097 ; n12098
g11843 and n11841_not n12098_not ; n12099
g11844 and n12095_not n12098_not ; n12100
g11845 and n12096_not n12100 ; n12101
g11846 and n12099_not n12101_not ; n12102
g11847 and b[44] n1302 ; n12103
g11848 and b[42] n1391 ; n12104
g11849 and b[43] n1297 ; n12105
g11850 and n12104_not n12105_not ; n12106
g11851 and n12103_not n12106 ; n12107
g11852 and n1305 n7072 ; n12108
g11853 and n12107 n12108_not ; n12109
g11854 and a[17] n12109_not ; n12110
g11855 and a[17] n12110_not ; n12111
g11856 and n12109_not n12110_not ; n12112
g11857 and n12111_not n12112_not ; n12113
g11858 and n12102_not n12113_not ; n12114
g11859 and n12102_not n12114_not ; n12115
g11860 and n12113_not n12114_not ; n12116
g11861 and n12115_not n12116_not ; n12117
g11862 and n11768_not n12117 ; n12118
g11863 and n11768 n12117_not ; n12119
g11864 and n12118_not n12119_not ; n12120
g11865 and b[47] n951 ; n12121
g11866 and b[45] n1056 ; n12122
g11867 and b[46] n946 ; n12123
g11868 and n12122_not n12123_not ; n12124
g11869 and n12121_not n12124 ; n12125
g11870 and n954 n7703 ; n12126
g11871 and n12125 n12126_not ; n12127
g11872 and a[14] n12127_not ; n12128
g11873 and a[14] n12128_not ; n12129
g11874 and n12127_not n12128_not ; n12130
g11875 and n12129_not n12130_not ; n12131
g11876 and n12120_not n12131_not ; n12132
g11877 and n12120 n12131 ; n12133
g11878 and n12132_not n12133_not ; n12134
g11879 and n11840_not n12134 ; n12135
g11880 and n11840 n12134_not ; n12136
g11881 and n12135_not n12136_not ; n12137
g11882 and n11839_not n12137 ; n12138
g11883 and n12137 n12138_not ; n12139
g11884 and n11839_not n12138_not ; n12140
g11885 and n12139_not n12140_not ; n12141
g11886 and n11828_not n12141_not ; n12142
g11887 and n11828 n12141 ; n12143
g11888 and n12142_not n12143_not ; n12144
g11889 and n11827_not n12144 ; n12145
g11890 and n11827_not n12145_not ; n12146
g11891 and n12144 n12145_not ; n12147
g11892 and n12146_not n12147_not ; n12148
g11893 and n11816_not n12148_not ; n12149
g11894 and n11816_not n12149_not ; n12150
g11895 and n12148_not n12149_not ; n12151
g11896 and n12150_not n12151_not ; n12152
g11897 and b[56] n362 ; n12153
g11898 and b[54] n403 ; n12154
g11899 and b[55] n357 ; n12155
g11900 and n12154_not n12155_not ; n12156
g11901 and n12153_not n12156 ; n12157
g11902 and n365 n10708 ; n12158
g11903 and n12157 n12158_not ; n12159
g11904 and a[5] n12159_not ; n12160
g11905 and a[5] n12160_not ; n12161
g11906 and n12159_not n12160_not ; n12162
g11907 and n12161_not n12162_not ; n12163
g11908 and n12152_not n12163_not ; n12164
g11909 and n12152_not n12164_not ; n12165
g11910 and n12163_not n12164_not ; n12166
g11911 and n12165_not n12166_not ; n12167
g11912 and b[59] n266 ; n12168
g11913 and b[57] n284 ; n12169
g11914 and b[58] n261 ; n12170
g11915 and n12169_not n12170_not ; n12171
g11916 and n12168_not n12171 ; n12172
g11917 and n11432_not n11434_not ; n12173
g11918 and b[58]_not b[59]_not ; n12174
g11919 and b[58] b[59] ; n12175
g11920 and n12174_not n12175_not ; n12176
g11921 and n12173_not n12176 ; n12177
g11922 and n12173 n12176_not ; n12178
g11923 and n12177_not n12178_not ; n12179
g11924 and n269 n12179 ; n12180
g11925 and n12172 n12180_not ; n12181
g11926 and a[2] n12181_not ; n12182
g11927 and a[2] n12182_not ; n12183
g11928 and n12181_not n12182_not ; n12184
g11929 and n12183_not n12184_not ; n12185
g11930 and n12167_not n12185 ; n12186
g11931 and n12167 n12185_not ; n12187
g11932 and n12186_not n12187_not ; n12188
g11933 and n11815_not n12188_not ; n12189
g11934 and n11815_not n12189_not ; n12190
g11935 and n12188_not n12189_not ; n12191
g11936 and n12190_not n12191_not ; n12192
g11937 and n11814_not n12192_not ; n12193
g11938 and n11814 n12191_not ; n12194
g11939 and n12190_not n12194 ; n12195
g11940 and n12193_not n12195_not ; f[59]
g11941 and n12189_not n12193_not ; n12197
g11942 and n12167_not n12185_not ; n12198
g11943 and n12164_not n12198_not ; n12199
g11944 and b[60] n266 ; n12200
g11945 and b[58] n284 ; n12201
g11946 and b[59] n261 ; n12202
g11947 and n12201_not n12202_not ; n12203
g11948 and n12200_not n12203 ; n12204
g11949 and n12175_not n12177_not ; n12205
g11950 and b[59]_not b[60]_not ; n12206
g11951 and b[59] b[60] ; n12207
g11952 and n12206_not n12207_not ; n12208
g11953 and n12205_not n12208 ; n12209
g11954 and n12205 n12208_not ; n12210
g11955 and n12209_not n12210_not ; n12211
g11956 and n269 n12211 ; n12212
g11957 and n12204 n12212_not ; n12213
g11958 and a[2] n12213_not ; n12214
g11959 and a[2] n12214_not ; n12215
g11960 and n12213_not n12214_not ; n12216
g11961 and n12215_not n12216_not ; n12217
g11962 and b[57] n362 ; n12218
g11963 and b[55] n403 ; n12219
g11964 and b[56] n357 ; n12220
g11965 and n12219_not n12220_not ; n12221
g11966 and n12218_not n12221 ; n12222
g11967 and n365 n11410 ; n12223
g11968 and n12222 n12223_not ; n12224
g11969 and a[5] n12224_not ; n12225
g11970 and a[5] n12225_not ; n12226
g11971 and n12224_not n12225_not ; n12227
g11972 and n12226_not n12227_not ; n12228
g11973 and n12145_not n12149_not ; n12229
g11974 and b[54] n511 ; n12230
g11975 and b[52] n541 ; n12231
g11976 and b[53] n506 ; n12232
g11977 and n12231_not n12232_not ; n12233
g11978 and n12230_not n12233 ; n12234
g11979 and n514 n9998 ; n12235
g11980 and n12234 n12235_not ; n12236
g11981 and a[8] n12236_not ; n12237
g11982 and a[8] n12237_not ; n12238
g11983 and n12236_not n12237_not ; n12239
g11984 and n12238_not n12239_not ; n12240
g11985 and n12138_not n12142_not ; n12241
g11986 and b[51] n700 ; n12242
g11987 and b[49] n767 ; n12243
g11988 and b[50] n695 ; n12244
g11989 and n12243_not n12244_not ; n12245
g11990 and n12242_not n12245 ; n12246
g11991 and n703 n8976 ; n12247
g11992 and n12246 n12247_not ; n12248
g11993 and a[11] n12248_not ; n12249
g11994 and a[11] n12249_not ; n12250
g11995 and n12248_not n12249_not ; n12251
g11996 and n12250_not n12251_not ; n12252
g11997 and n12132_not n12135_not ; n12253
g11998 and b[48] n951 ; n12254
g11999 and b[46] n1056 ; n12255
g12000 and b[47] n946 ; n12256
g12001 and n12255_not n12256_not ; n12257
g12002 and n12254_not n12257 ; n12258
g12003 and n954 n8009 ; n12259
g12004 and n12258 n12259_not ; n12260
g12005 and a[14] n12260_not ; n12261
g12006 and a[14] n12261_not ; n12262
g12007 and n12260_not n12261_not ; n12263
g12008 and n12262_not n12263_not ; n12264
g12009 and n11768_not n12117_not ; n12265
g12010 and n12114_not n12265_not ; n12266
g12011 and b[45] n1302 ; n12267
g12012 and b[43] n1391 ; n12268
g12013 and b[44] n1297 ; n12269
g12014 and n12268_not n12269_not ; n12270
g12015 and n12267_not n12270 ; n12271
g12016 and n1305 n7361 ; n12272
g12017 and n12271 n12272_not ; n12273
g12018 and a[17] n12273_not ; n12274
g12019 and a[17] n12274_not ; n12275
g12020 and n12273_not n12274_not ; n12276
g12021 and n12275_not n12276_not ; n12277
g12022 and n12057_not n12063_not ; n12278
g12023 and n12052_not n12054_not ; n12279
g12024 and b[33] n3050 ; n12280
g12025 and b[31] n3243 ; n12281
g12026 and b[32] n3045 ; n12282
g12027 and n12281_not n12282_not ; n12283
g12028 and n12280_not n12283 ; n12284
g12029 and n3053 n4223 ; n12285
g12030 and n12284 n12285_not ; n12286
g12031 and a[29] n12286_not ; n12287
g12032 and a[29] n12287_not ; n12288
g12033 and n12286_not n12287_not ; n12289
g12034 and n12288_not n12289_not ; n12290
g12035 and n11618_not n11981_not ; n12291
g12036 and n11978_not n12291_not ; n12292
g12037 and b[21] n5777 ; n12293
g12038 and b[19] n6059 ; n12294
g12039 and b[20] n5772 ; n12295
g12040 and n12294_not n12295_not ; n12296
g12041 and n12293_not n12296 ; n12297
g12042 and n1984 n5780 ; n12298
g12043 and n12297 n12298_not ; n12299
g12044 and a[41] n12299_not ; n12300
g12045 and a[41] n12300_not ; n12301
g12046 and n12299_not n12300_not ; n12302
g12047 and n12301_not n12302_not ; n12303
g12048 and n11959_not n11963_not ; n12304
g12049 and b[18] n6595 ; n12305
g12050 and b[16] n6902 ; n12306
g12051 and b[17] n6590 ; n12307
g12052 and n12306_not n12307_not ; n12308
g12053 and n12305_not n12308 ; n12309
g12054 and n1566 n6598 ; n12310
g12055 and n12309 n12310_not ; n12311
g12056 and a[44] n12311_not ; n12312
g12057 and a[44] n12312_not ; n12313
g12058 and n12311_not n12312_not ; n12314
g12059 and n12313_not n12314_not ; n12315
g12060 and n11952_not n11956_not ; n12316
g12061 and b[15] n7446 ; n12317
g12062 and b[13] n7787 ; n12318
g12063 and b[14] n7441 ; n12319
g12064 and n12318_not n12319_not ; n12320
g12065 and n12317_not n12320 ; n12321
g12066 and n1131 n7449 ; n12322
g12067 and n12321 n12322_not ; n12323
g12068 and a[47] n12323_not ; n12324
g12069 and a[47] n12324_not ; n12325
g12070 and n12323_not n12324_not ; n12326
g12071 and n12325_not n12326_not ; n12327
g12072 and n11947_not n11949_not ; n12328
g12073 and b[12] n8362 ; n12329
g12074 and b[10] n8715 ; n12330
g12075 and b[11] n8357 ; n12331
g12076 and n12330_not n12331_not ; n12332
g12077 and n12329_not n12332 ; n12333
g12078 and n842 n8365 ; n12334
g12079 and n12333 n12334_not ; n12335
g12080 and a[50] n12335_not ; n12336
g12081 and a[50] n12336_not ; n12337
g12082 and n12335_not n12336_not ; n12338
g12083 and n12337_not n12338_not ; n12339
g12084 and n11941_not n11943_not ; n12340
g12085 and b[6] n10426 ; n12341
g12086 and b[4] n10796 ; n12342
g12087 and b[5] n10421 ; n12343
g12088 and n12342_not n12343_not ; n12344
g12089 and n12341_not n12344 ; n12345
g12090 and n459 n10429 ; n12346
g12091 and n12345 n12346_not ; n12347
g12092 and a[56] n12347_not ; n12348
g12093 and a[56] n12348_not ; n12349
g12094 and n12347_not n12348_not ; n12350
g12095 and n12349_not n12350_not ; n12351
g12096 and a[59] a[60]_not ; n12352
g12097 and a[59]_not a[60] ; n12353
g12098 and n12352_not n12353_not ; n12354
g12099 and b[0] n12354_not ; n12355
g12100 and n11908_not n12355 ; n12356
g12101 and n11908 n12355_not ; n12357
g12102 and n12356_not n12357_not ; n12358
g12103 and b[3] n11531 ; n12359
g12104 and b[1] n11896 ; n12360
g12105 and b[2] n11526 ; n12361
g12106 and n12360_not n12361_not ; n12362
g12107 and n12359_not n12362 ; n12363
g12108 and n318 n11534 ; n12364
g12109 and n12363 n12364_not ; n12365
g12110 and a[59] n12365_not ; n12366
g12111 and a[59] n12366_not ; n12367
g12112 and n12365_not n12366_not ; n12368
g12113 and n12367_not n12368_not ; n12369
g12114 and n12358_not n12369_not ; n12370
g12115 and n12358 n12369 ; n12371
g12116 and n12370_not n12371_not ; n12372
g12117 and n12351_not n12372 ; n12373
g12118 and n12372 n12373_not ; n12374
g12119 and n12351_not n12373_not ; n12375
g12120 and n12374_not n12375_not ; n12376
g12121 and n11926_not n12376 ; n12377
g12122 and n11926 n12376_not ; n12378
g12123 and n12377_not n12378_not ; n12379
g12124 and b[9] n9339 ; n12380
g12125 and b[7] n9732 ; n12381
g12126 and b[8] n9334 ; n12382
g12127 and n12381_not n12382_not ; n12383
g12128 and n12380_not n12383 ; n12384
g12129 and n651 n9342 ; n12385
g12130 and n12384 n12385_not ; n12386
g12131 and a[53] n12386_not ; n12387
g12132 and a[53] n12387_not ; n12388
g12133 and n12386_not n12387_not ; n12389
g12134 and n12388_not n12389_not ; n12390
g12135 and n12379_not n12390_not ; n12391
g12136 and n12379 n12390 ; n12392
g12137 and n12391_not n12392_not ; n12393
g12138 and n12340_not n12393 ; n12394
g12139 and n12340 n12393_not ; n12395
g12140 and n12394_not n12395_not ; n12396
g12141 and n12339 n12396_not ; n12397
g12142 and n12339_not n12396 ; n12398
g12143 and n12397_not n12398_not ; n12399
g12144 and n12328_not n12399 ; n12400
g12145 and n12328 n12399_not ; n12401
g12146 and n12400_not n12401_not ; n12402
g12147 and n12327_not n12402 ; n12403
g12148 and n12327 n12402_not ; n12404
g12149 and n12403_not n12404_not ; n12405
g12150 and n12316_not n12405 ; n12406
g12151 and n12316 n12405_not ; n12407
g12152 and n12406_not n12407_not ; n12408
g12153 and n12315_not n12408 ; n12409
g12154 and n12315_not n12409_not ; n12410
g12155 and n12408 n12409_not ; n12411
g12156 and n12410_not n12411_not ; n12412
g12157 and n12304_not n12412_not ; n12413
g12158 and n12304 n12411_not ; n12414
g12159 and n12410_not n12414 ; n12415
g12160 and n12413_not n12415_not ; n12416
g12161 and n12303_not n12416 ; n12417
g12162 and n12303 n12416_not ; n12418
g12163 and n12417_not n12418_not ; n12419
g12164 and n12292_not n12419 ; n12420
g12165 and n12292 n12419_not ; n12421
g12166 and n12420_not n12421_not ; n12422
g12167 and b[24] n5035 ; n12423
g12168 and b[22] n5277 ; n12424
g12169 and b[23] n5030 ; n12425
g12170 and n12424_not n12425_not ; n12426
g12171 and n12423_not n12426 ; n12427
g12172 and n2458 n5038 ; n12428
g12173 and n12427 n12428_not ; n12429
g12174 and a[38] n12429_not ; n12430
g12175 and a[38] n12430_not ; n12431
g12176 and n12429_not n12430_not ; n12432
g12177 and n12431_not n12432_not ; n12433
g12178 and n12422 n12433_not ; n12434
g12179 and n12422 n12434_not ; n12435
g12180 and n12433_not n12434_not ; n12436
g12181 and n12435_not n12436_not ; n12437
g12182 and n11996_not n12000_not ; n12438
g12183 and n12437 n12438 ; n12439
g12184 and n12437_not n12438_not ; n12440
g12185 and n12439_not n12440_not ; n12441
g12186 and b[27] n4287 ; n12442
g12187 and b[25] n4532 ; n12443
g12188 and b[26] n4282 ; n12444
g12189 and n12443_not n12444_not ; n12445
g12190 and n12442_not n12445 ; n12446
g12191 and n2990 n4290 ; n12447
g12192 and n12446 n12447_not ; n12448
g12193 and a[35] n12448_not ; n12449
g12194 and a[35] n12449_not ; n12450
g12195 and n12448_not n12449_not ; n12451
g12196 and n12450_not n12451_not ; n12452
g12197 and n12441 n12452_not ; n12453
g12198 and n12441 n12453_not ; n12454
g12199 and n12452_not n12453_not ; n12455
g12200 and n12454_not n12455_not ; n12456
g12201 and n12013_not n12019_not ; n12457
g12202 and n12456 n12457 ; n12458
g12203 and n12456_not n12457_not ; n12459
g12204 and n12458_not n12459_not ; n12460
g12205 and b[30] n3638 ; n12461
g12206 and b[28] n3843 ; n12462
g12207 and b[29] n3633 ; n12463
g12208 and n12462_not n12463_not ; n12464
g12209 and n12461_not n12464 ; n12465
g12210 and n3577 n3641 ; n12466
g12211 and n12465 n12466_not ; n12467
g12212 and a[32] n12467_not ; n12468
g12213 and a[32] n12468_not ; n12469
g12214 and n12467_not n12468_not ; n12470
g12215 and n12469_not n12470_not ; n12471
g12216 and n12460_not n12471 ; n12472
g12217 and n12460 n12471_not ; n12473
g12218 and n12472_not n12473_not ; n12474
g12219 and n12037_not n12474 ; n12475
g12220 and n12037 n12474_not ; n12476
g12221 and n12475_not n12476_not ; n12477
g12222 and n12290_not n12477 ; n12478
g12223 and n12477 n12478_not ; n12479
g12224 and n12290_not n12478_not ; n12480
g12225 and n12479_not n12480_not ; n12481
g12226 and n12279_not n12481 ; n12482
g12227 and n12279 n12481_not ; n12483
g12228 and n12482_not n12483_not ; n12484
g12229 and b[36] n2539 ; n12485
g12230 and b[34] n2685 ; n12486
g12231 and b[35] n2534 ; n12487
g12232 and n12486_not n12487_not ; n12488
g12233 and n12485_not n12488 ; n12489
g12234 and n2542 n4922 ; n12490
g12235 and n12489 n12490_not ; n12491
g12236 and a[26] n12491_not ; n12492
g12237 and a[26] n12492_not ; n12493
g12238 and n12491_not n12492_not ; n12494
g12239 and n12493_not n12494_not ; n12495
g12240 and n12484_not n12495_not ; n12496
g12241 and n12484 n12495 ; n12497
g12242 and n12496_not n12497_not ; n12498
g12243 and n12278 n12498_not ; n12499
g12244 and n12278_not n12498 ; n12500
g12245 and n12499_not n12500_not ; n12501
g12246 and b[39] n2048 ; n12502
g12247 and b[37] n2198 ; n12503
g12248 and b[38] n2043 ; n12504
g12249 and n12503_not n12504_not ; n12505
g12250 and n12502_not n12505 ; n12506
g12251 and n2051 n5451 ; n12507
g12252 and n12506 n12507_not ; n12508
g12253 and a[23] n12508_not ; n12509
g12254 and a[23] n12509_not ; n12510
g12255 and n12508_not n12509_not ; n12511
g12256 and n12510_not n12511_not ; n12512
g12257 and n12501 n12512_not ; n12513
g12258 and n12501 n12513_not ; n12514
g12259 and n12512_not n12513_not ; n12515
g12260 and n12514_not n12515_not ; n12516
g12261 and n12076_not n12082_not ; n12517
g12262 and n12516 n12517 ; n12518
g12263 and n12516_not n12517_not ; n12519
g12264 and n12518_not n12519_not ; n12520
g12265 and b[42] n1627 ; n12521
g12266 and b[40] n1763 ; n12522
g12267 and b[41] n1622 ; n12523
g12268 and n12522_not n12523_not ; n12524
g12269 and n12521_not n12524 ; n12525
g12270 and n1630 n6489 ; n12526
g12271 and n12525 n12526_not ; n12527
g12272 and a[20] n12527_not ; n12528
g12273 and a[20] n12528_not ; n12529
g12274 and n12527_not n12528_not ; n12530
g12275 and n12529_not n12530_not ; n12531
g12276 and n12520_not n12531 ; n12532
g12277 and n12520 n12531_not ; n12533
g12278 and n12532_not n12533_not ; n12534
g12279 and n12100_not n12534 ; n12535
g12280 and n12100 n12534_not ; n12536
g12281 and n12535_not n12536_not ; n12537
g12282 and n12277_not n12537 ; n12538
g12283 and n12277_not n12538_not ; n12539
g12284 and n12537 n12538_not ; n12540
g12285 and n12539_not n12540_not ; n12541
g12286 and n12266_not n12541_not ; n12542
g12287 and n12266 n12540_not ; n12543
g12288 and n12539_not n12543 ; n12544
g12289 and n12542_not n12544_not ; n12545
g12290 and n12264_not n12545 ; n12546
g12291 and n12264_not n12546_not ; n12547
g12292 and n12545 n12546_not ; n12548
g12293 and n12547_not n12548_not ; n12549
g12294 and n12253_not n12549_not ; n12550
g12295 and n12253 n12548_not ; n12551
g12296 and n12547_not n12551 ; n12552
g12297 and n12550_not n12552_not ; n12553
g12298 and n12252_not n12553 ; n12554
g12299 and n12252_not n12554_not ; n12555
g12300 and n12553 n12554_not ; n12556
g12301 and n12555_not n12556_not ; n12557
g12302 and n12241_not n12557_not ; n12558
g12303 and n12241 n12556_not ; n12559
g12304 and n12555_not n12559 ; n12560
g12305 and n12558_not n12560_not ; n12561
g12306 and n12240_not n12561 ; n12562
g12307 and n12240 n12561_not ; n12563
g12308 and n12562_not n12563_not ; n12564
g12309 and n12229_not n12564 ; n12565
g12310 and n12229 n12564_not ; n12566
g12311 and n12565_not n12566_not ; n12567
g12312 and n12228_not n12567 ; n12568
g12313 and n12228 n12567_not ; n12569
g12314 and n12568_not n12569_not ; n12570
g12315 and n12217_not n12570 ; n12571
g12316 and n12217 n12570_not ; n12572
g12317 and n12571_not n12572_not ; n12573
g12318 and n12199_not n12573 ; n12574
g12319 and n12199 n12573_not ; n12575
g12320 and n12574_not n12575_not ; n12576
g12321 and n12197_not n12576 ; n12577
g12322 and n12197 n12576_not ; n12578
g12323 and n12577_not n12578_not ; f[60]
g12324 and b[55] n511 ; n12580
g12325 and b[53] n541 ; n12581
g12326 and b[54] n506 ; n12582
g12327 and n12581_not n12582_not ; n12583
g12328 and n12580_not n12583 ; n12584
g12329 and n514 n10684 ; n12585
g12330 and n12584 n12585_not ; n12586
g12331 and a[8] n12586_not ; n12587
g12332 and a[8] n12587_not ; n12588
g12333 and n12586_not n12587_not ; n12589
g12334 and n12588_not n12589_not ; n12590
g12335 and n12554_not n12558_not ; n12591
g12336 and b[52] n700 ; n12592
g12337 and b[50] n767 ; n12593
g12338 and b[51] n695 ; n12594
g12339 and n12593_not n12594_not ; n12595
g12340 and n12592_not n12595 ; n12596
g12341 and n703 n9628 ; n12597
g12342 and n12596 n12597_not ; n12598
g12343 and a[11] n12598_not ; n12599
g12344 and a[11] n12599_not ; n12600
g12345 and n12598_not n12599_not ; n12601
g12346 and n12600_not n12601_not ; n12602
g12347 and n12546_not n12550_not ; n12603
g12348 and b[49] n951 ; n12604
g12349 and b[47] n1056 ; n12605
g12350 and b[48] n946 ; n12606
g12351 and n12605_not n12606_not ; n12607
g12352 and n12604_not n12607 ; n12608
g12353 and n954 n8625 ; n12609
g12354 and n12608 n12609_not ; n12610
g12355 and a[14] n12610_not ; n12611
g12356 and a[14] n12611_not ; n12612
g12357 and n12610_not n12611_not ; n12613
g12358 and n12612_not n12613_not ; n12614
g12359 and n12538_not n12542_not ; n12615
g12360 and n12533_not n12535_not ; n12616
g12361 and n12279_not n12481_not ; n12617
g12362 and n12478_not n12617_not ; n12618
g12363 and n12473_not n12475_not ; n12619
g12364 and n12409_not n12413_not ; n12620
g12365 and n12398_not n12400_not ; n12621
g12366 and b[10] n9339 ; n12622
g12367 and b[8] n9732 ; n12623
g12368 and b[9] n9334 ; n12624
g12369 and n12623_not n12624_not ; n12625
g12370 and n12622_not n12625 ; n12626
g12371 and n738 n9342 ; n12627
g12372 and n12626 n12627_not ; n12628
g12373 and a[53] n12628_not ; n12629
g12374 and a[53] n12629_not ; n12630
g12375 and n12628_not n12629_not ; n12631
g12376 and n12630_not n12631_not ; n12632
g12377 and n11926_not n12376_not ; n12633
g12378 and n12373_not n12633_not ; n12634
g12379 and b[7] n10426 ; n12635
g12380 and b[5] n10796 ; n12636
g12381 and b[6] n10421 ; n12637
g12382 and n12636_not n12637_not ; n12638
g12383 and n12635_not n12638 ; n12639
g12384 and n484 n10429 ; n12640
g12385 and n12639 n12640_not ; n12641
g12386 and a[56] n12641_not ; n12642
g12387 and a[56] n12642_not ; n12643
g12388 and n12641_not n12642_not ; n12644
g12389 and n12643_not n12644_not ; n12645
g12390 and n11908 n12355 ; n12646
g12391 and n12370_not n12646_not ; n12647
g12392 and b[4] n11531 ; n12648
g12393 and b[2] n11896 ; n12649
g12394 and b[3] n11526 ; n12650
g12395 and n12649_not n12650_not ; n12651
g12396 and n12648_not n12651 ; n12652
g12397 and n346 n11534 ; n12653
g12398 and n12652 n12653_not ; n12654
g12399 and a[59] n12654_not ; n12655
g12400 and a[59] n12655_not ; n12656
g12401 and n12654_not n12655_not ; n12657
g12402 and n12656_not n12657_not ; n12658
g12403 and a[62] n12355_not ; n12659
g12404 and a[60]_not a[61] ; n12660
g12405 and a[60] a[61]_not ; n12661
g12406 and n12660_not n12661_not ; n12662
g12407 and n12354 n12662_not ; n12663
g12408 and b[0] n12663 ; n12664
g12409 and a[61]_not a[62] ; n12665
g12410 and a[61] a[62]_not ; n12666
g12411 and n12665_not n12666_not ; n12667
g12412 and n12354_not n12667 ; n12668
g12413 and b[1] n12668 ; n12669
g12414 and n12664_not n12669_not ; n12670
g12415 and n12354_not n12667_not ; n12671
g12416 and n272_not n12671 ; n12672
g12417 and n12670 n12672_not ; n12673
g12418 and a[62] n12673_not ; n12674
g12419 and a[62] n12674_not ; n12675
g12420 and n12673_not n12674_not ; n12676
g12421 and n12675_not n12676_not ; n12677
g12422 and n12659 n12677_not ; n12678
g12423 and n12659_not n12677 ; n12679
g12424 and n12678_not n12679_not ; n12680
g12425 and n12658 n12680_not ; n12681
g12426 and n12658_not n12680 ; n12682
g12427 and n12681_not n12682_not ; n12683
g12428 and n12647_not n12683 ; n12684
g12429 and n12647 n12683_not ; n12685
g12430 and n12684_not n12685_not ; n12686
g12431 and n12645 n12686_not ; n12687
g12432 and n12645_not n12686 ; n12688
g12433 and n12687_not n12688_not ; n12689
g12434 and n12634_not n12689 ; n12690
g12435 and n12634 n12689_not ; n12691
g12436 and n12690_not n12691_not ; n12692
g12437 and n12632_not n12692 ; n12693
g12438 and n12692 n12693_not ; n12694
g12439 and n12632_not n12693_not ; n12695
g12440 and n12694_not n12695_not ; n12696
g12441 and n12391_not n12394_not ; n12697
g12442 and n12696 n12697 ; n12698
g12443 and n12696_not n12697_not ; n12699
g12444 and n12698_not n12699_not ; n12700
g12445 and b[13] n8362 ; n12701
g12446 and b[11] n8715 ; n12702
g12447 and b[12] n8357 ; n12703
g12448 and n12702_not n12703_not ; n12704
g12449 and n12701_not n12704 ; n12705
g12450 and n1008 n8365 ; n12706
g12451 and n12705 n12706_not ; n12707
g12452 and a[50] n12707_not ; n12708
g12453 and a[50] n12708_not ; n12709
g12454 and n12707_not n12708_not ; n12710
g12455 and n12709_not n12710_not ; n12711
g12456 and n12700 n12711_not ; n12712
g12457 and n12700_not n12711 ; n12713
g12458 and n12621_not n12713_not ; n12714
g12459 and n12712_not n12714 ; n12715
g12460 and n12621_not n12715_not ; n12716
g12461 and n12712_not n12715_not ; n12717
g12462 and n12713_not n12717 ; n12718
g12463 and n12716_not n12718_not ; n12719
g12464 and b[16] n7446 ; n12720
g12465 and b[14] n7787 ; n12721
g12466 and b[15] n7441 ; n12722
g12467 and n12721_not n12722_not ; n12723
g12468 and n12720_not n12723 ; n12724
g12469 and n1237 n7449 ; n12725
g12470 and n12724 n12725_not ; n12726
g12471 and a[47] n12726_not ; n12727
g12472 and a[47] n12727_not ; n12728
g12473 and n12726_not n12727_not ; n12729
g12474 and n12728_not n12729_not ; n12730
g12475 and n12719_not n12730_not ; n12731
g12476 and n12719_not n12731_not ; n12732
g12477 and n12730_not n12731_not ; n12733
g12478 and n12732_not n12733_not ; n12734
g12479 and n12403_not n12406_not ; n12735
g12480 and n12734 n12735 ; n12736
g12481 and n12734_not n12735_not ; n12737
g12482 and n12736_not n12737_not ; n12738
g12483 and b[19] n6595 ; n12739
g12484 and b[17] n6902 ; n12740
g12485 and b[18] n6590 ; n12741
g12486 and n12740_not n12741_not ; n12742
g12487 and n12739_not n12742 ; n12743
g12488 and n1708 n6598 ; n12744
g12489 and n12743 n12744_not ; n12745
g12490 and a[44] n12745_not ; n12746
g12491 and a[44] n12746_not ; n12747
g12492 and n12745_not n12746_not ; n12748
g12493 and n12747_not n12748_not ; n12749
g12494 and n12738 n12749_not ; n12750
g12495 and n12738_not n12749 ; n12751
g12496 and n12620_not n12751_not ; n12752
g12497 and n12750_not n12752 ; n12753
g12498 and n12620_not n12753_not ; n12754
g12499 and n12750_not n12753_not ; n12755
g12500 and n12751_not n12755 ; n12756
g12501 and n12754_not n12756_not ; n12757
g12502 and b[22] n5777 ; n12758
g12503 and b[20] n6059 ; n12759
g12504 and b[21] n5772 ; n12760
g12505 and n12759_not n12760_not ; n12761
g12506 and n12758_not n12761 ; n12762
g12507 and n2145 n5780 ; n12763
g12508 and n12762 n12763_not ; n12764
g12509 and a[41] n12764_not ; n12765
g12510 and a[41] n12765_not ; n12766
g12511 and n12764_not n12765_not ; n12767
g12512 and n12766_not n12767_not ; n12768
g12513 and n12757_not n12768_not ; n12769
g12514 and n12757_not n12769_not ; n12770
g12515 and n12768_not n12769_not ; n12771
g12516 and n12770_not n12771_not ; n12772
g12517 and n12417_not n12420_not ; n12773
g12518 and n12772 n12773 ; n12774
g12519 and n12772_not n12773_not ; n12775
g12520 and n12774_not n12775_not ; n12776
g12521 and b[25] n5035 ; n12777
g12522 and b[23] n5277 ; n12778
g12523 and b[24] n5030 ; n12779
g12524 and n12778_not n12779_not ; n12780
g12525 and n12777_not n12780 ; n12781
g12526 and n2485 n5038 ; n12782
g12527 and n12781 n12782_not ; n12783
g12528 and a[38] n12783_not ; n12784
g12529 and a[38] n12784_not ; n12785
g12530 and n12783_not n12784_not ; n12786
g12531 and n12785_not n12786_not ; n12787
g12532 and n12776 n12787_not ; n12788
g12533 and n12776 n12788_not ; n12789
g12534 and n12787_not n12788_not ; n12790
g12535 and n12789_not n12790_not ; n12791
g12536 and n12434_not n12440_not ; n12792
g12537 and n12791 n12792 ; n12793
g12538 and n12791_not n12792_not ; n12794
g12539 and n12793_not n12794_not ; n12795
g12540 and b[28] n4287 ; n12796
g12541 and b[26] n4532 ; n12797
g12542 and b[27] n4282 ; n12798
g12543 and n12797_not n12798_not ; n12799
g12544 and n12796_not n12799 ; n12800
g12545 and n3189 n4290 ; n12801
g12546 and n12800 n12801_not ; n12802
g12547 and a[35] n12802_not ; n12803
g12548 and a[35] n12803_not ; n12804
g12549 and n12802_not n12803_not ; n12805
g12550 and n12804_not n12805_not ; n12806
g12551 and n12795 n12806_not ; n12807
g12552 and n12795 n12807_not ; n12808
g12553 and n12806_not n12807_not ; n12809
g12554 and n12808_not n12809_not ; n12810
g12555 and n12453_not n12459_not ; n12811
g12556 and n12810 n12811 ; n12812
g12557 and n12810_not n12811_not ; n12813
g12558 and n12812_not n12813_not ; n12814
g12559 and b[31] n3638 ; n12815
g12560 and b[29] n3843 ; n12816
g12561 and b[30] n3633 ; n12817
g12562 and n12816_not n12817_not ; n12818
g12563 and n12815_not n12818 ; n12819
g12564 and n3641 n3796 ; n12820
g12565 and n12819 n12820_not ; n12821
g12566 and a[32] n12821_not ; n12822
g12567 and a[32] n12822_not ; n12823
g12568 and n12821_not n12822_not ; n12824
g12569 and n12823_not n12824_not ; n12825
g12570 and n12814 n12825_not ; n12826
g12571 and n12814 n12826_not ; n12827
g12572 and n12825_not n12826_not ; n12828
g12573 and n12827_not n12828_not ; n12829
g12574 and n12619_not n12829 ; n12830
g12575 and n12619 n12829_not ; n12831
g12576 and n12830_not n12831_not ; n12832
g12577 and b[34] n3050 ; n12833
g12578 and b[32] n3243 ; n12834
g12579 and b[33] n3045 ; n12835
g12580 and n12834_not n12835_not ; n12836
g12581 and n12833_not n12836 ; n12837
g12582 and n3053 n4466 ; n12838
g12583 and n12837 n12838_not ; n12839
g12584 and a[29] n12839_not ; n12840
g12585 and a[29] n12840_not ; n12841
g12586 and n12839_not n12840_not ; n12842
g12587 and n12841_not n12842_not ; n12843
g12588 and n12832_not n12843_not ; n12844
g12589 and n12832 n12843 ; n12845
g12590 and n12844_not n12845_not ; n12846
g12591 and n12618 n12846_not ; n12847
g12592 and n12618_not n12846 ; n12848
g12593 and n12847_not n12848_not ; n12849
g12594 and b[37] n2539 ; n12850
g12595 and b[35] n2685 ; n12851
g12596 and b[36] n2534 ; n12852
g12597 and n12851_not n12852_not ; n12853
g12598 and n12850_not n12853 ; n12854
g12599 and n2542 n5181 ; n12855
g12600 and n12854 n12855_not ; n12856
g12601 and a[26] n12856_not ; n12857
g12602 and a[26] n12857_not ; n12858
g12603 and n12856_not n12857_not ; n12859
g12604 and n12858_not n12859_not ; n12860
g12605 and n12849 n12860_not ; n12861
g12606 and n12849 n12861_not ; n12862
g12607 and n12860_not n12861_not ; n12863
g12608 and n12862_not n12863_not ; n12864
g12609 and n12496_not n12500_not ; n12865
g12610 and n12864 n12865 ; n12866
g12611 and n12864_not n12865_not ; n12867
g12612 and n12866_not n12867_not ; n12868
g12613 and b[40] n2048 ; n12869
g12614 and b[38] n2198 ; n12870
g12615 and b[39] n2043 ; n12871
g12616 and n12870_not n12871_not ; n12872
g12617 and n12869_not n12872 ; n12873
g12618 and n2051 n5955 ; n12874
g12619 and n12873 n12874_not ; n12875
g12620 and a[23] n12875_not ; n12876
g12621 and a[23] n12876_not ; n12877
g12622 and n12875_not n12876_not ; n12878
g12623 and n12877_not n12878_not ; n12879
g12624 and n12868 n12879_not ; n12880
g12625 and n12868 n12880_not ; n12881
g12626 and n12879_not n12880_not ; n12882
g12627 and n12881_not n12882_not ; n12883
g12628 and n12513_not n12519_not ; n12884
g12629 and n12883 n12884 ; n12885
g12630 and n12883_not n12884_not ; n12886
g12631 and n12885_not n12886_not ; n12887
g12632 and b[43] n1627 ; n12888
g12633 and b[41] n1763 ; n12889
g12634 and b[42] n1622 ; n12890
g12635 and n12889_not n12890_not ; n12891
g12636 and n12888_not n12891 ; n12892
g12637 and n1630 n6515 ; n12893
g12638 and n12892 n12893_not ; n12894
g12639 and a[20] n12894_not ; n12895
g12640 and a[20] n12895_not ; n12896
g12641 and n12894_not n12895_not ; n12897
g12642 and n12896_not n12897_not ; n12898
g12643 and n12887 n12898_not ; n12899
g12644 and n12887_not n12898 ; n12900
g12645 and n12616_not n12900_not ; n12901
g12646 and n12899_not n12901 ; n12902
g12647 and n12616_not n12902_not ; n12903
g12648 and n12899_not n12902_not ; n12904
g12649 and n12900_not n12904 ; n12905
g12650 and n12903_not n12905_not ; n12906
g12651 and b[46] n1302 ; n12907
g12652 and b[44] n1391 ; n12908
g12653 and b[45] n1297 ; n12909
g12654 and n12908_not n12909_not ; n12910
g12655 and n12907_not n12910 ; n12911
g12656 and n1305 n7677 ; n12912
g12657 and n12911 n12912_not ; n12913
g12658 and a[17] n12913_not ; n12914
g12659 and a[17] n12914_not ; n12915
g12660 and n12913_not n12914_not ; n12916
g12661 and n12915_not n12916_not ; n12917
g12662 and n12906 n12917 ; n12918
g12663 and n12906_not n12917_not ; n12919
g12664 and n12918_not n12919_not ; n12920
g12665 and n12615_not n12920 ; n12921
g12666 and n12615 n12920_not ; n12922
g12667 and n12921_not n12922_not ; n12923
g12668 and n12614 n12923_not ; n12924
g12669 and n12614_not n12923 ; n12925
g12670 and n12924_not n12925_not ; n12926
g12671 and n12603_not n12926 ; n12927
g12672 and n12603 n12926_not ; n12928
g12673 and n12927_not n12928_not ; n12929
g12674 and n12602 n12929_not ; n12930
g12675 and n12602_not n12929 ; n12931
g12676 and n12930_not n12931_not ; n12932
g12677 and n12591_not n12932 ; n12933
g12678 and n12591 n12932_not ; n12934
g12679 and n12933_not n12934_not ; n12935
g12680 and n12590_not n12935 ; n12936
g12681 and n12935 n12936_not ; n12937
g12682 and n12590_not n12936_not ; n12938
g12683 and n12937_not n12938_not ; n12939
g12684 and n12562_not n12565_not ; n12940
g12685 and n12939 n12940 ; n12941
g12686 and n12939_not n12940_not ; n12942
g12687 and n12941_not n12942_not ; n12943
g12688 and b[58] n362 ; n12944
g12689 and b[56] n403 ; n12945
g12690 and b[57] n357 ; n12946
g12691 and n12945_not n12946_not ; n12947
g12692 and n12944_not n12947 ; n12948
g12693 and n365 n11436 ; n12949
g12694 and n12948 n12949_not ; n12950
g12695 and a[5] n12950_not ; n12951
g12696 and a[5] n12951_not ; n12952
g12697 and n12950_not n12951_not ; n12953
g12698 and n12952_not n12953_not ; n12954
g12699 and n12943_not n12954 ; n12955
g12700 and n12943 n12954_not ; n12956
g12701 and n12955_not n12956_not ; n12957
g12702 and b[61] n266 ; n12958
g12703 and b[59] n284 ; n12959
g12704 and b[60] n261 ; n12960
g12705 and n12959_not n12960_not ; n12961
g12706 and n12958_not n12961 ; n12962
g12707 and n12207_not n12209_not ; n12963
g12708 and b[60]_not b[61]_not ; n12964
g12709 and b[60] b[61] ; n12965
g12710 and n12964_not n12965_not ; n12966
g12711 and n12963_not n12966 ; n12967
g12712 and n12963 n12966_not ; n12968
g12713 and n12967_not n12968_not ; n12969
g12714 and n269 n12969 ; n12970
g12715 and n12962 n12970_not ; n12971
g12716 and a[2] n12971_not ; n12972
g12717 and a[2] n12972_not ; n12973
g12718 and n12971_not n12972_not ; n12974
g12719 and n12973_not n12974_not ; n12975
g12720 and n12957 n12975_not ; n12976
g12721 and n12957 n12976_not ; n12977
g12722 and n12975_not n12976_not ; n12978
g12723 and n12977_not n12978_not ; n12979
g12724 and n12568_not n12571_not ; n12980
g12725 and n12979 n12980 ; n12981
g12726 and n12979_not n12980_not ; n12982
g12727 and n12981_not n12982_not ; n12983
g12728 and n12574_not n12577_not ; n12984
g12729 and n12983 n12984_not ; n12985
g12730 and n12983_not n12984 ; n12986
g12731 and n12985_not n12986_not ; f[61]
g12732 and n12982_not n12985_not ; n12988
g12733 and n12956_not n12976_not ; n12989
g12734 and n12931_not n12933_not ; n12990
g12735 and n12925_not n12927_not ; n12991
g12736 and b[50] n951 ; n12992
g12737 and b[48] n1056 ; n12993
g12738 and b[49] n946 ; n12994
g12739 and n12993_not n12994_not ; n12995
g12740 and n12992_not n12995 ; n12996
g12741 and n954 n8949 ; n12997
g12742 and n12996 n12997_not ; n12998
g12743 and a[14] n12998_not ; n12999
g12744 and a[14] n12999_not ; n13000
g12745 and n12998_not n12999_not ; n13001
g12746 and n13000_not n13001_not ; n13002
g12747 and n12919_not n12921_not ; n13003
g12748 and n12880_not n12886_not ; n13004
g12749 and n12619_not n12829_not ; n13005
g12750 and n12826_not n13005_not ; n13006
g12751 and n12769_not n12775_not ; n13007
g12752 and n12731_not n12737_not ; n13008
g12753 and b[17] n7446 ; n13009
g12754 and b[15] n7787 ; n13010
g12755 and b[16] n7441 ; n13011
g12756 and n13010_not n13011_not ; n13012
g12757 and n13009_not n13012 ; n13013
g12758 and n1356 n7449 ; n13014
g12759 and n13013 n13014_not ; n13015
g12760 and a[47] n13015_not ; n13016
g12761 and a[47] n13016_not ; n13017
g12762 and n13015_not n13016_not ; n13018
g12763 and n13017_not n13018_not ; n13019
g12764 and b[14] n8362 ; n13020
g12765 and b[12] n8715 ; n13021
g12766 and b[13] n8357 ; n13022
g12767 and n13021_not n13022_not ; n13023
g12768 and n13020_not n13023 ; n13024
g12769 and n1034 n8365 ; n13025
g12770 and n13024 n13025_not ; n13026
g12771 and a[50] n13026_not ; n13027
g12772 and a[50] n13027_not ; n13028
g12773 and n13026_not n13027_not ; n13029
g12774 and n13028_not n13029_not ; n13030
g12775 and n12693_not n12699_not ; n13031
g12776 and b[11] n9339 ; n13032
g12777 and b[9] n9732 ; n13033
g12778 and b[10] n9334 ; n13034
g12779 and n13033_not n13034_not ; n13035
g12780 and n13032_not n13035 ; n13036
g12781 and n818 n9342 ; n13037
g12782 and n13036 n13037_not ; n13038
g12783 and a[53] n13038_not ; n13039
g12784 and a[53] n13039_not ; n13040
g12785 and n13038_not n13039_not ; n13041
g12786 and n13040_not n13041_not ; n13042
g12787 and n12688_not n12690_not ; n13043
g12788 and n12682_not n12684_not ; n13044
g12789 and b[2] n12668 ; n13045
g12790 and n12354 n12667_not ; n13046
g12791 and n12662 n13046 ; n13047
g12792 and b[0] n13047 ; n13048
g12793 and b[1] n12663 ; n13049
g12794 and n13048_not n13049_not ; n13050
g12795 and n13045_not n13050 ; n13051
g12796 and n296 n12671 ; n13052
g12797 and n13051 n13052_not ; n13053
g12798 and a[62] n13053_not ; n13054
g12799 and a[62] n13054_not ; n13055
g12800 and n13053_not n13054_not ; n13056
g12801 and n13055_not n13056_not ; n13057
g12802 and n12678_not n13057 ; n13058
g12803 and n12678 n13057_not ; n13059
g12804 and n13058_not n13059_not ; n13060
g12805 and b[5] n11531 ; n13061
g12806 and b[3] n11896 ; n13062
g12807 and b[4] n11526 ; n13063
g12808 and n13062_not n13063_not ; n13064
g12809 and n13061_not n13064 ; n13065
g12810 and n394 n11534 ; n13066
g12811 and n13065 n13066_not ; n13067
g12812 and a[59] n13067_not ; n13068
g12813 and a[59] n13068_not ; n13069
g12814 and n13067_not n13068_not ; n13070
g12815 and n13069_not n13070_not ; n13071
g12816 and n13060 n13071_not ; n13072
g12817 and n13060_not n13071 ; n13073
g12818 and n13044_not n13073_not ; n13074
g12819 and n13072_not n13074 ; n13075
g12820 and n13044_not n13075_not ; n13076
g12821 and n13072_not n13075_not ; n13077
g12822 and n13073_not n13077 ; n13078
g12823 and n13076_not n13078_not ; n13079
g12824 and b[8] n10426 ; n13080
g12825 and b[6] n10796 ; n13081
g12826 and b[7] n10421 ; n13082
g12827 and n13081_not n13082_not ; n13083
g12828 and n13080_not n13083 ; n13084
g12829 and n585 n10429 ; n13085
g12830 and n13084 n13085_not ; n13086
g12831 and a[56] n13086_not ; n13087
g12832 and a[56] n13087_not ; n13088
g12833 and n13086_not n13087_not ; n13089
g12834 and n13088_not n13089_not ; n13090
g12835 and n13079 n13090 ; n13091
g12836 and n13079_not n13090_not ; n13092
g12837 and n13091_not n13092_not ; n13093
g12838 and n13043_not n13093 ; n13094
g12839 and n13043 n13093_not ; n13095
g12840 and n13094_not n13095_not ; n13096
g12841 and n13042 n13096_not ; n13097
g12842 and n13042_not n13096 ; n13098
g12843 and n13097_not n13098_not ; n13099
g12844 and n13031_not n13099 ; n13100
g12845 and n13031 n13099_not ; n13101
g12846 and n13100_not n13101_not ; n13102
g12847 and n13030_not n13102 ; n13103
g12848 and n13102 n13103_not ; n13104
g12849 and n13030_not n13103_not ; n13105
g12850 and n13104_not n13105_not ; n13106
g12851 and n12717_not n13106_not ; n13107
g12852 and n12717 n13106 ; n13108
g12853 and n13107_not n13108_not ; n13109
g12854 and n13019_not n13109 ; n13110
g12855 and n13019_not n13110_not ; n13111
g12856 and n13109 n13110_not ; n13112
g12857 and n13111_not n13112_not ; n13113
g12858 and n13008_not n13113_not ; n13114
g12859 and n13008_not n13114_not ; n13115
g12860 and n13113_not n13114_not ; n13116
g12861 and n13115_not n13116_not ; n13117
g12862 and b[20] n6595 ; n13118
g12863 and b[18] n6902 ; n13119
g12864 and b[19] n6590 ; n13120
g12865 and n13119_not n13120_not ; n13121
g12866 and n13118_not n13121 ; n13122
g12867 and n1846 n6598 ; n13123
g12868 and n13122 n13123_not ; n13124
g12869 and a[44] n13124_not ; n13125
g12870 and a[44] n13125_not ; n13126
g12871 and n13124_not n13125_not ; n13127
g12872 and n13126_not n13127_not ; n13128
g12873 and n13117_not n13128_not ; n13129
g12874 and n13117_not n13129_not ; n13130
g12875 and n13128_not n13129_not ; n13131
g12876 and n13130_not n13131_not ; n13132
g12877 and n12755_not n13132 ; n13133
g12878 and n12755 n13132_not ; n13134
g12879 and n13133_not n13134_not ; n13135
g12880 and b[23] n5777 ; n13136
g12881 and b[21] n6059 ; n13137
g12882 and b[22] n5772 ; n13138
g12883 and n13137_not n13138_not ; n13139
g12884 and n13136_not n13139 ; n13140
g12885 and n2300 n5780 ; n13141
g12886 and n13140 n13141_not ; n13142
g12887 and a[41] n13142_not ; n13143
g12888 and a[41] n13143_not ; n13144
g12889 and n13142_not n13143_not ; n13145
g12890 and n13144_not n13145_not ; n13146
g12891 and n13135_not n13146_not ; n13147
g12892 and n13135 n13146 ; n13148
g12893 and n13147_not n13148_not ; n13149
g12894 and n13007 n13149_not ; n13150
g12895 and n13007_not n13149 ; n13151
g12896 and n13150_not n13151_not ; n13152
g12897 and b[26] n5035 ; n13153
g12898 and b[24] n5277 ; n13154
g12899 and b[25] n5030 ; n13155
g12900 and n13154_not n13155_not ; n13156
g12901 and n13153_not n13156 ; n13157
g12902 and n2813 n5038 ; n13158
g12903 and n13157 n13158_not ; n13159
g12904 and a[38] n13159_not ; n13160
g12905 and a[38] n13160_not ; n13161
g12906 and n13159_not n13160_not ; n13162
g12907 and n13161_not n13162_not ; n13163
g12908 and n13152 n13163_not ; n13164
g12909 and n13152 n13164_not ; n13165
g12910 and n13163_not n13164_not ; n13166
g12911 and n13165_not n13166_not ; n13167
g12912 and n12788_not n12794_not ; n13168
g12913 and n13167 n13168 ; n13169
g12914 and n13167_not n13168_not ; n13170
g12915 and n13169_not n13170_not ; n13171
g12916 and b[29] n4287 ; n13172
g12917 and b[27] n4532 ; n13173
g12918 and b[28] n4282 ; n13174
g12919 and n13173_not n13174_not ; n13175
g12920 and n13172_not n13175 ; n13176
g12921 and n3383 n4290 ; n13177
g12922 and n13176 n13177_not ; n13178
g12923 and a[35] n13178_not ; n13179
g12924 and a[35] n13179_not ; n13180
g12925 and n13178_not n13179_not ; n13181
g12926 and n13180_not n13181_not ; n13182
g12927 and n13171 n13182_not ; n13183
g12928 and n13171 n13183_not ; n13184
g12929 and n13182_not n13183_not ; n13185
g12930 and n13184_not n13185_not ; n13186
g12931 and n12807_not n12813_not ; n13187
g12932 and n13186 n13187 ; n13188
g12933 and n13186_not n13187_not ; n13189
g12934 and n13188_not n13189_not ; n13190
g12935 and b[32] n3638 ; n13191
g12936 and b[30] n3843 ; n13192
g12937 and b[31] n3633 ; n13193
g12938 and n13192_not n13193_not ; n13194
g12939 and n13191_not n13194 ; n13195
g12940 and n3641 n4013 ; n13196
g12941 and n13195 n13196_not ; n13197
g12942 and a[32] n13197_not ; n13198
g12943 and a[32] n13198_not ; n13199
g12944 and n13197_not n13198_not ; n13200
g12945 and n13199_not n13200_not ; n13201
g12946 and n13190 n13201_not ; n13202
g12947 and n13190_not n13201 ; n13203
g12948 and n13006_not n13203_not ; n13204
g12949 and n13202_not n13204 ; n13205
g12950 and n13006_not n13205_not ; n13206
g12951 and n13202_not n13205_not ; n13207
g12952 and n13203_not n13207 ; n13208
g12953 and n13206_not n13208_not ; n13209
g12954 and b[35] n3050 ; n13210
g12955 and b[33] n3243 ; n13211
g12956 and b[34] n3045 ; n13212
g12957 and n13211_not n13212_not ; n13213
g12958 and n13210_not n13213 ; n13214
g12959 and n3053 n4696 ; n13215
g12960 and n13214 n13215_not ; n13216
g12961 and a[29] n13216_not ; n13217
g12962 and a[29] n13217_not ; n13218
g12963 and n13216_not n13217_not ; n13219
g12964 and n13218_not n13219_not ; n13220
g12965 and n13209_not n13220_not ; n13221
g12966 and n13209_not n13221_not ; n13222
g12967 and n13220_not n13221_not ; n13223
g12968 and n13222_not n13223_not ; n13224
g12969 and n12844_not n12848_not ; n13225
g12970 and n13224 n13225 ; n13226
g12971 and n13224_not n13225_not ; n13227
g12972 and n13226_not n13227_not ; n13228
g12973 and b[38] n2539 ; n13229
g12974 and b[36] n2685 ; n13230
g12975 and b[37] n2534 ; n13231
g12976 and n13230_not n13231_not ; n13232
g12977 and n13229_not n13232 ; n13233
g12978 and n2542 n5205 ; n13234
g12979 and n13233 n13234_not ; n13235
g12980 and a[26] n13235_not ; n13236
g12981 and a[26] n13236_not ; n13237
g12982 and n13235_not n13236_not ; n13238
g12983 and n13237_not n13238_not ; n13239
g12984 and n13228 n13239_not ; n13240
g12985 and n13228 n13240_not ; n13241
g12986 and n13239_not n13240_not ; n13242
g12987 and n13241_not n13242_not ; n13243
g12988 and n12861_not n12867_not ; n13244
g12989 and n13243 n13244 ; n13245
g12990 and n13243_not n13244_not ; n13246
g12991 and n13245_not n13246_not ; n13247
g12992 and b[41] n2048 ; n13248
g12993 and b[39] n2198 ; n13249
g12994 and b[40] n2043 ; n13250
g12995 and n13249_not n13250_not ; n13251
g12996 and n13248_not n13251 ; n13252
g12997 and n2051 n6219 ; n13253
g12998 and n13252 n13253_not ; n13254
g12999 and a[23] n13254_not ; n13255
g13000 and a[23] n13255_not ; n13256
g13001 and n13254_not n13255_not ; n13257
g13002 and n13256_not n13257_not ; n13258
g13003 and n13247 n13258_not ; n13259
g13004 and n13247_not n13258 ; n13260
g13005 and n13004_not n13260_not ; n13261
g13006 and n13259_not n13261 ; n13262
g13007 and n13004_not n13262_not ; n13263
g13008 and n13259_not n13262_not ; n13264
g13009 and n13260_not n13264 ; n13265
g13010 and n13263_not n13265_not ; n13266
g13011 and b[44] n1627 ; n13267
g13012 and b[42] n1763 ; n13268
g13013 and b[43] n1622 ; n13269
g13014 and n13268_not n13269_not ; n13270
g13015 and n13267_not n13270 ; n13271
g13016 and n1630 n7072 ; n13272
g13017 and n13271 n13272_not ; n13273
g13018 and a[20] n13273_not ; n13274
g13019 and a[20] n13274_not ; n13275
g13020 and n13273_not n13274_not ; n13276
g13021 and n13275_not n13276_not ; n13277
g13022 and n13266_not n13277_not ; n13278
g13023 and n13266_not n13278_not ; n13279
g13024 and n13277_not n13278_not ; n13280
g13025 and n13279_not n13280_not ; n13281
g13026 and n12904_not n13281 ; n13282
g13027 and n12904 n13281_not ; n13283
g13028 and n13282_not n13283_not ; n13284
g13029 and b[47] n1302 ; n13285
g13030 and b[45] n1391 ; n13286
g13031 and b[46] n1297 ; n13287
g13032 and n13286_not n13287_not ; n13288
g13033 and n13285_not n13288 ; n13289
g13034 and n1305 n7703 ; n13290
g13035 and n13289 n13290_not ; n13291
g13036 and a[17] n13291_not ; n13292
g13037 and a[17] n13292_not ; n13293
g13038 and n13291_not n13292_not ; n13294
g13039 and n13293_not n13294_not ; n13295
g13040 and n13284_not n13295_not ; n13296
g13041 and n13284 n13295 ; n13297
g13042 and n13296_not n13297_not ; n13298
g13043 and n13003_not n13298 ; n13299
g13044 and n13003 n13298_not ; n13300
g13045 and n13299_not n13300_not ; n13301
g13046 and n13002_not n13301 ; n13302
g13047 and n13301 n13302_not ; n13303
g13048 and n13002_not n13302_not ; n13304
g13049 and n13303_not n13304_not ; n13305
g13050 and n12991_not n13305 ; n13306
g13051 and n12991 n13305_not ; n13307
g13052 and n13306_not n13307_not ; n13308
g13053 and b[53] n700 ; n13309
g13054 and b[51] n767 ; n13310
g13055 and b[52] n695 ; n13311
g13056 and n13310_not n13311_not ; n13312
g13057 and n13309_not n13312 ; n13313
g13058 and n703 n9972 ; n13314
g13059 and n13313 n13314_not ; n13315
g13060 and a[11] n13315_not ; n13316
g13061 and a[11] n13316_not ; n13317
g13062 and n13315_not n13316_not ; n13318
g13063 and n13317_not n13318_not ; n13319
g13064 and n13308_not n13319_not ; n13320
g13065 and n13308 n13319 ; n13321
g13066 and n13320_not n13321_not ; n13322
g13067 and n12990_not n13322 ; n13323
g13068 and n12990 n13322_not ; n13324
g13069 and n13323_not n13324_not ; n13325
g13070 and b[56] n511 ; n13326
g13071 and b[54] n541 ; n13327
g13072 and b[55] n506 ; n13328
g13073 and n13327_not n13328_not ; n13329
g13074 and n13326_not n13329 ; n13330
g13075 and n514 n10708 ; n13331
g13076 and n13330 n13331_not ; n13332
g13077 and a[8] n13332_not ; n13333
g13078 and a[8] n13333_not ; n13334
g13079 and n13332_not n13333_not ; n13335
g13080 and n13334_not n13335_not ; n13336
g13081 and n13325_not n13336 ; n13337
g13082 and n13325 n13336_not ; n13338
g13083 and n13337_not n13338_not ; n13339
g13084 and b[59] n362 ; n13340
g13085 and b[57] n403 ; n13341
g13086 and b[58] n357 ; n13342
g13087 and n13341_not n13342_not ; n13343
g13088 and n13340_not n13343 ; n13344
g13089 and n365 n12179 ; n13345
g13090 and n13344 n13345_not ; n13346
g13091 and a[5] n13346_not ; n13347
g13092 and a[5] n13347_not ; n13348
g13093 and n13346_not n13347_not ; n13349
g13094 and n13348_not n13349_not ; n13350
g13095 and n13339 n13350_not ; n13351
g13096 and n13339 n13351_not ; n13352
g13097 and n13350_not n13351_not ; n13353
g13098 and n13352_not n13353_not ; n13354
g13099 and n12936_not n12942_not ; n13355
g13100 and n13354 n13355 ; n13356
g13101 and n13354_not n13355_not ; n13357
g13102 and n13356_not n13357_not ; n13358
g13103 and b[62] n266 ; n13359
g13104 and b[60] n284 ; n13360
g13105 and b[61] n261 ; n13361
g13106 and n13360_not n13361_not ; n13362
g13107 and n13359_not n13362 ; n13363
g13108 and n12965_not n12967_not ; n13364
g13109 and b[61]_not b[62]_not ; n13365
g13110 and b[61] b[62] ; n13366
g13111 and n13365_not n13366_not ; n13367
g13112 and n13364_not n13367 ; n13368
g13113 and n13364 n13367_not ; n13369
g13114 and n13368_not n13369_not ; n13370
g13115 and n269 n13370 ; n13371
g13116 and n13363 n13371_not ; n13372
g13117 and a[2] n13372_not ; n13373
g13118 and a[2] n13373_not ; n13374
g13119 and n13372_not n13373_not ; n13375
g13120 and n13374_not n13375_not ; n13376
g13121 and n13358_not n13376 ; n13377
g13122 and n13358 n13376_not ; n13378
g13123 and n13377_not n13378_not ; n13379
g13124 and n12989_not n13379 ; n13380
g13125 and n12989 n13379_not ; n13381
g13126 and n13380_not n13381_not ; n13382
g13127 and n12988_not n13382 ; n13383
g13128 and n12988 n13382_not ; n13384
g13129 and n13383_not n13384_not ; f[62]
g13130 and n12991_not n13305_not ; n13386
g13131 and n13302_not n13386_not ; n13387
g13132 and b[51] n951 ; n13388
g13133 and b[49] n1056 ; n13389
g13134 and b[50] n946 ; n13390
g13135 and n13389_not n13390_not ; n13391
g13136 and n13388_not n13391 ; n13392
g13137 and n954 n8976 ; n13393
g13138 and n13392 n13393_not ; n13394
g13139 and a[14] n13394_not ; n13395
g13140 and a[14] n13395_not ; n13396
g13141 and n13394_not n13395_not ; n13397
g13142 and n13396_not n13397_not ; n13398
g13143 and n13296_not n13299_not ; n13399
g13144 and b[48] n1302 ; n13400
g13145 and b[46] n1391 ; n13401
g13146 and b[47] n1297 ; n13402
g13147 and n13401_not n13402_not ; n13403
g13148 and n13400_not n13403 ; n13404
g13149 and n1305 n8009 ; n13405
g13150 and n13404 n13405_not ; n13406
g13151 and a[17] n13406_not ; n13407
g13152 and a[17] n13407_not ; n13408
g13153 and n13406_not n13407_not ; n13409
g13154 and n13408_not n13409_not ; n13410
g13155 and n12904_not n13281_not ; n13411
g13156 and n13278_not n13411_not ; n13412
g13157 and b[45] n1627 ; n13413
g13158 and b[43] n1763 ; n13414
g13159 and b[44] n1622 ; n13415
g13160 and n13414_not n13415_not ; n13416
g13161 and n13413_not n13416 ; n13417
g13162 and n1630 n7361 ; n13418
g13163 and n13417 n13418_not ; n13419
g13164 and a[20] n13419_not ; n13420
g13165 and a[20] n13420_not ; n13421
g13166 and n13419_not n13420_not ; n13422
g13167 and n13421_not n13422_not ; n13423
g13168 and b[42] n2048 ; n13424
g13169 and b[40] n2198 ; n13425
g13170 and b[41] n2043 ; n13426
g13171 and n13425_not n13426_not ; n13427
g13172 and n13424_not n13427 ; n13428
g13173 and n2051 n6489 ; n13429
g13174 and n13428 n13429_not ; n13430
g13175 and a[23] n13430_not ; n13431
g13176 and a[23] n13431_not ; n13432
g13177 and n13430_not n13431_not ; n13433
g13178 and n13432_not n13433_not ; n13434
g13179 and n13240_not n13246_not ; n13435
g13180 and n13221_not n13227_not ; n13436
g13181 and b[33] n3638 ; n13437
g13182 and b[31] n3843 ; n13438
g13183 and b[32] n3633 ; n13439
g13184 and n13438_not n13439_not ; n13440
g13185 and n13437_not n13440 ; n13441
g13186 and n3641 n4223 ; n13442
g13187 and n13441 n13442_not ; n13443
g13188 and a[32] n13443_not ; n13444
g13189 and a[32] n13444_not ; n13445
g13190 and n13443_not n13444_not ; n13446
g13191 and n13445_not n13446_not ; n13447
g13192 and n12755_not n13132_not ; n13448
g13193 and n13129_not n13448_not ; n13449
g13194 and b[21] n6595 ; n13450
g13195 and b[19] n6902 ; n13451
g13196 and b[20] n6590 ; n13452
g13197 and n13451_not n13452_not ; n13453
g13198 and n13450_not n13453 ; n13454
g13199 and n1984 n6598 ; n13455
g13200 and n13454 n13455_not ; n13456
g13201 and a[44] n13456_not ; n13457
g13202 and a[44] n13457_not ; n13458
g13203 and n13456_not n13457_not ; n13459
g13204 and n13458_not n13459_not ; n13460
g13205 and n13110_not n13114_not ; n13461
g13206 and b[15] n8362 ; n13462
g13207 and b[13] n8715 ; n13463
g13208 and b[14] n8357 ; n13464
g13209 and n13463_not n13464_not ; n13465
g13210 and n13462_not n13465 ; n13466
g13211 and n1131 n8365 ; n13467
g13212 and n13466 n13467_not ; n13468
g13213 and a[50] n13468_not ; n13469
g13214 and a[50] n13469_not ; n13470
g13215 and n13468_not n13469_not ; n13471
g13216 and n13470_not n13471_not ; n13472
g13217 and n13098_not n13100_not ; n13473
g13218 and n13092_not n13094_not ; n13474
g13219 and b[9] n10426 ; n13475
g13220 and b[7] n10796 ; n13476
g13221 and b[8] n10421 ; n13477
g13222 and n13476_not n13477_not ; n13478
g13223 and n13475_not n13478 ; n13479
g13224 and n651 n10429 ; n13480
g13225 and n13479 n13480_not ; n13481
g13226 and a[56] n13481_not ; n13482
g13227 and a[56] n13482_not ; n13483
g13228 and n13481_not n13482_not ; n13484
g13229 and n13483_not n13484_not ; n13485
g13230 and a[62] a[63]_not ; n13486
g13231 and a[62]_not a[63] ; n13487
g13232 and n13486_not n13487_not ; n13488
g13233 and b[0] n13488_not ; n13489
g13234 and n13059 n13489 ; n13490
g13235 and n13059 n13490_not ; n13491
g13236 and n13489 n13490_not ; n13492
g13237 and n13491_not n13492_not ; n13493
g13238 and b[3] n12668 ; n13494
g13239 and b[1] n13047 ; n13495
g13240 and b[2] n12663 ; n13496
g13241 and n13495_not n13496_not ; n13497
g13242 and n13494_not n13497 ; n13498
g13243 and n318 n12671 ; n13499
g13244 and n13498 n13499_not ; n13500
g13245 and a[62] n13500_not ; n13501
g13246 and a[62] n13501_not ; n13502
g13247 and n13500_not n13501_not ; n13503
g13248 and n13502_not n13503_not ; n13504
g13249 and n13493_not n13504_not ; n13505
g13250 and n13493_not n13505_not ; n13506
g13251 and n13504_not n13505_not ; n13507
g13252 and n13506_not n13507_not ; n13508
g13253 and b[6] n11531 ; n13509
g13254 and b[4] n11896 ; n13510
g13255 and b[5] n11526 ; n13511
g13256 and n13510_not n13511_not ; n13512
g13257 and n13509_not n13512 ; n13513
g13258 and n459 n11534 ; n13514
g13259 and n13513 n13514_not ; n13515
g13260 and a[59] n13515_not ; n13516
g13261 and a[59] n13516_not ; n13517
g13262 and n13515_not n13516_not ; n13518
g13263 and n13517_not n13518_not ; n13519
g13264 and n13508 n13519 ; n13520
g13265 and n13508_not n13519_not ; n13521
g13266 and n13520_not n13521_not ; n13522
g13267 and n13077_not n13522 ; n13523
g13268 and n13077 n13522_not ; n13524
g13269 and n13523_not n13524_not ; n13525
g13270 and n13485_not n13525 ; n13526
g13271 and n13525 n13526_not ; n13527
g13272 and n13485_not n13526_not ; n13528
g13273 and n13527_not n13528_not ; n13529
g13274 and n13474_not n13529 ; n13530
g13275 and n13474 n13529_not ; n13531
g13276 and n13530_not n13531_not ; n13532
g13277 and b[12] n9339 ; n13533
g13278 and b[10] n9732 ; n13534
g13279 and b[11] n9334 ; n13535
g13280 and n13534_not n13535_not ; n13536
g13281 and n13533_not n13536 ; n13537
g13282 and n842 n9342 ; n13538
g13283 and n13537 n13538_not ; n13539
g13284 and a[53] n13539_not ; n13540
g13285 and a[53] n13540_not ; n13541
g13286 and n13539_not n13540_not ; n13542
g13287 and n13541_not n13542_not ; n13543
g13288 and n13532 n13543 ; n13544
g13289 and n13532_not n13543_not ; n13545
g13290 and n13544_not n13545_not ; n13546
g13291 and n13473_not n13546 ; n13547
g13292 and n13473 n13546_not ; n13548
g13293 and n13547_not n13548_not ; n13549
g13294 and n13472_not n13549 ; n13550
g13295 and n13549 n13550_not ; n13551
g13296 and n13472_not n13550_not ; n13552
g13297 and n13551_not n13552_not ; n13553
g13298 and n13103_not n13107_not ; n13554
g13299 and n13553 n13554 ; n13555
g13300 and n13553_not n13554_not ; n13556
g13301 and n13555_not n13556_not ; n13557
g13302 and b[18] n7446 ; n13558
g13303 and b[16] n7787 ; n13559
g13304 and b[17] n7441 ; n13560
g13305 and n13559_not n13560_not ; n13561
g13306 and n13558_not n13561 ; n13562
g13307 and n1566 n7449 ; n13563
g13308 and n13562 n13563_not ; n13564
g13309 and a[47] n13564_not ; n13565
g13310 and a[47] n13565_not ; n13566
g13311 and n13564_not n13565_not ; n13567
g13312 and n13566_not n13567_not ; n13568
g13313 and n13557_not n13568 ; n13569
g13314 and n13557 n13568_not ; n13570
g13315 and n13569_not n13570_not ; n13571
g13316 and n13461_not n13571 ; n13572
g13317 and n13461 n13571_not ; n13573
g13318 and n13572_not n13573_not ; n13574
g13319 and n13460_not n13574 ; n13575
g13320 and n13460 n13574_not ; n13576
g13321 and n13575_not n13576_not ; n13577
g13322 and n13449_not n13577 ; n13578
g13323 and n13449 n13577_not ; n13579
g13324 and n13578_not n13579_not ; n13580
g13325 and b[24] n5777 ; n13581
g13326 and b[22] n6059 ; n13582
g13327 and b[23] n5772 ; n13583
g13328 and n13582_not n13583_not ; n13584
g13329 and n13581_not n13584 ; n13585
g13330 and n2458 n5780 ; n13586
g13331 and n13585 n13586_not ; n13587
g13332 and a[41] n13587_not ; n13588
g13333 and a[41] n13588_not ; n13589
g13334 and n13587_not n13588_not ; n13590
g13335 and n13589_not n13590_not ; n13591
g13336 and n13580 n13591_not ; n13592
g13337 and n13580 n13592_not ; n13593
g13338 and n13591_not n13592_not ; n13594
g13339 and n13593_not n13594_not ; n13595
g13340 and n13147_not n13151_not ; n13596
g13341 and n13595 n13596 ; n13597
g13342 and n13595_not n13596_not ; n13598
g13343 and n13597_not n13598_not ; n13599
g13344 and b[27] n5035 ; n13600
g13345 and b[25] n5277 ; n13601
g13346 and b[26] n5030 ; n13602
g13347 and n13601_not n13602_not ; n13603
g13348 and n13600_not n13603 ; n13604
g13349 and n2990 n5038 ; n13605
g13350 and n13604 n13605_not ; n13606
g13351 and a[38] n13606_not ; n13607
g13352 and a[38] n13607_not ; n13608
g13353 and n13606_not n13607_not ; n13609
g13354 and n13608_not n13609_not ; n13610
g13355 and n13599 n13610_not ; n13611
g13356 and n13599 n13611_not ; n13612
g13357 and n13610_not n13611_not ; n13613
g13358 and n13612_not n13613_not ; n13614
g13359 and n13164_not n13170_not ; n13615
g13360 and n13614 n13615 ; n13616
g13361 and n13614_not n13615_not ; n13617
g13362 and n13616_not n13617_not ; n13618
g13363 and b[30] n4287 ; n13619
g13364 and b[28] n4532 ; n13620
g13365 and b[29] n4282 ; n13621
g13366 and n13620_not n13621_not ; n13622
g13367 and n13619_not n13622 ; n13623
g13368 and n3577 n4290 ; n13624
g13369 and n13623 n13624_not ; n13625
g13370 and a[35] n13625_not ; n13626
g13371 and a[35] n13626_not ; n13627
g13372 and n13625_not n13626_not ; n13628
g13373 and n13627_not n13628_not ; n13629
g13374 and n13618_not n13629 ; n13630
g13375 and n13618 n13629_not ; n13631
g13376 and n13630_not n13631_not ; n13632
g13377 and n13183_not n13189_not ; n13633
g13378 and n13632 n13633_not ; n13634
g13379 and n13632_not n13633 ; n13635
g13380 and n13634_not n13635_not ; n13636
g13381 and n13447_not n13636 ; n13637
g13382 and n13636 n13637_not ; n13638
g13383 and n13447_not n13637_not ; n13639
g13384 and n13638_not n13639_not ; n13640
g13385 and n13207_not n13640 ; n13641
g13386 and n13207 n13640_not ; n13642
g13387 and n13641_not n13642_not ; n13643
g13388 and b[36] n3050 ; n13644
g13389 and b[34] n3243 ; n13645
g13390 and b[35] n3045 ; n13646
g13391 and n13645_not n13646_not ; n13647
g13392 and n13644_not n13647 ; n13648
g13393 and n3053 n4922 ; n13649
g13394 and n13648 n13649_not ; n13650
g13395 and a[29] n13650_not ; n13651
g13396 and a[29] n13651_not ; n13652
g13397 and n13650_not n13651_not ; n13653
g13398 and n13652_not n13653_not ; n13654
g13399 and n13643_not n13654_not ; n13655
g13400 and n13643 n13654 ; n13656
g13401 and n13655_not n13656_not ; n13657
g13402 and n13436 n13657_not ; n13658
g13403 and n13436_not n13657 ; n13659
g13404 and n13658_not n13659_not ; n13660
g13405 and b[39] n2539 ; n13661
g13406 and b[37] n2685 ; n13662
g13407 and b[38] n2534 ; n13663
g13408 and n13662_not n13663_not ; n13664
g13409 and n13661_not n13664 ; n13665
g13410 and n2542 n5451 ; n13666
g13411 and n13665 n13666_not ; n13667
g13412 and a[26] n13667_not ; n13668
g13413 and a[26] n13668_not ; n13669
g13414 and n13667_not n13668_not ; n13670
g13415 and n13669_not n13670_not ; n13671
g13416 and n13660_not n13671 ; n13672
g13417 and n13660 n13671_not ; n13673
g13418 and n13672_not n13673_not ; n13674
g13419 and n13435_not n13674 ; n13675
g13420 and n13435 n13674_not ; n13676
g13421 and n13675_not n13676_not ; n13677
g13422 and n13434_not n13677 ; n13678
g13423 and n13434_not n13678_not ; n13679
g13424 and n13677 n13678_not ; n13680
g13425 and n13679_not n13680_not ; n13681
g13426 and n13264_not n13681_not ; n13682
g13427 and n13264 n13680_not ; n13683
g13428 and n13679_not n13683 ; n13684
g13429 and n13682_not n13684_not ; n13685
g13430 and n13423_not n13685 ; n13686
g13431 and n13423_not n13686_not ; n13687
g13432 and n13685 n13686_not ; n13688
g13433 and n13687_not n13688_not ; n13689
g13434 and n13412_not n13689_not ; n13690
g13435 and n13412 n13688_not ; n13691
g13436 and n13687_not n13691 ; n13692
g13437 and n13690_not n13692_not ; n13693
g13438 and n13410_not n13693 ; n13694
g13439 and n13410_not n13694_not ; n13695
g13440 and n13693 n13694_not ; n13696
g13441 and n13695_not n13696_not ; n13697
g13442 and n13399_not n13697_not ; n13698
g13443 and n13399 n13696_not ; n13699
g13444 and n13695_not n13699 ; n13700
g13445 and n13698_not n13700_not ; n13701
g13446 and n13398_not n13701 ; n13702
g13447 and n13398 n13701_not ; n13703
g13448 and n13702_not n13703_not ; n13704
g13449 and n13387_not n13704 ; n13705
g13450 and n13387 n13704_not ; n13706
g13451 and n13705_not n13706_not ; n13707
g13452 and b[54] n700 ; n13708
g13453 and b[52] n767 ; n13709
g13454 and b[53] n695 ; n13710
g13455 and n13709_not n13710_not ; n13711
g13456 and n13708_not n13711 ; n13712
g13457 and n703 n9998 ; n13713
g13458 and n13712 n13713_not ; n13714
g13459 and a[11] n13714_not ; n13715
g13460 and a[11] n13715_not ; n13716
g13461 and n13714_not n13715_not ; n13717
g13462 and n13716_not n13717_not ; n13718
g13463 and n13707 n13718_not ; n13719
g13464 and n13707 n13719_not ; n13720
g13465 and n13718_not n13719_not ; n13721
g13466 and n13720_not n13721_not ; n13722
g13467 and n13320_not n13323_not ; n13723
g13468 and n13722 n13723 ; n13724
g13469 and n13722_not n13723_not ; n13725
g13470 and n13724_not n13725_not ; n13726
g13471 and b[57] n511 ; n13727
g13472 and b[55] n541 ; n13728
g13473 and b[56] n506 ; n13729
g13474 and n13728_not n13729_not ; n13730
g13475 and n13727_not n13730 ; n13731
g13476 and n514 n11410 ; n13732
g13477 and n13731 n13732_not ; n13733
g13478 and a[8] n13733_not ; n13734
g13479 and a[8] n13734_not ; n13735
g13480 and n13733_not n13734_not ; n13736
g13481 and n13735_not n13736_not ; n13737
g13482 and n13726 n13737_not ; n13738
g13483 and n13726 n13738_not ; n13739
g13484 and n13737_not n13738_not ; n13740
g13485 and n13739_not n13740_not ; n13741
g13486 and b[60] n362 ; n13742
g13487 and b[58] n403 ; n13743
g13488 and b[59] n357 ; n13744
g13489 and n13743_not n13744_not ; n13745
g13490 and n13742_not n13745 ; n13746
g13491 and n365 n12211 ; n13747
g13492 and n13746 n13747_not ; n13748
g13493 and a[5] n13748_not ; n13749
g13494 and a[5] n13749_not ; n13750
g13495 and n13748_not n13749_not ; n13751
g13496 and n13750_not n13751_not ; n13752
g13497 and n13741_not n13752 ; n13753
g13498 and n13741 n13752_not ; n13754
g13499 and n13753_not n13754_not ; n13755
g13500 and n13338_not n13351_not ; n13756
g13501 and n13755 n13756 ; n13757
g13502 and n13755_not n13756_not ; n13758
g13503 and n13757_not n13758_not ; n13759
g13504 and b[63] n266 ; n13760
g13505 and b[61] n284 ; n13761
g13506 and b[62] n261 ; n13762
g13507 and n13761_not n13762_not ; n13763
g13508 and n13760_not n13763 ; n13764
g13509 and n13366_not n13368_not ; n13765
g13510 and b[62] b[63]_not ; n13766
g13511 and b[62]_not b[63] ; n13767
g13512 and n13766_not n13767_not ; n13768
g13513 and n13765_not n13768_not ; n13769
g13514 and n13765 n13768 ; n13770
g13515 and n13769_not n13770_not ; n13771
g13516 and n269 n13771 ; n13772
g13517 and n13764 n13772_not ; n13773
g13518 and a[2] n13773_not ; n13774
g13519 and a[2] n13774_not ; n13775
g13520 and n13773_not n13774_not ; n13776
g13521 and n13775_not n13776_not ; n13777
g13522 and n13759 n13777_not ; n13778
g13523 and n13759 n13778_not ; n13779
g13524 and n13777_not n13778_not ; n13780
g13525 and n13779_not n13780_not ; n13781
g13526 and n13357_not n13378_not ; n13782
g13527 and n13781_not n13782_not ; n13783
g13528 and n13781_not n13783_not ; n13784
g13529 and n13782_not n13783_not ; n13785
g13530 and n13784_not n13785_not ; n13786
g13531 and n13380_not n13383_not ; n13787
g13532 and n13786_not n13787_not ; n13788
g13533 and n13786 n13787 ; n13789
g13534 and n13788_not n13789_not ; f[63]
g13535 and n13783_not n13788_not ; n13791
g13536 and n13758_not n13778_not ; n13792
g13537 and b[62] n284 ; n13793
g13538 and b[63] n261 ; n13794
g13539 and n13793_not n13794_not ; n13795
g13540 and b[62]_not n13769_not ; n13796
g13541 and b[63] n13796_not ; n13797
g13542 and b[63] n13797_not ; n13798
g13543 and n13765_not n13766 ; n13799
g13544 and n13798_not n13799_not ; n13800
g13545 and n269 n13800_not ; n13801
g13546 and n13795 n13801_not ; n13802
g13547 and a[2] n13802_not ; n13803
g13548 and a[2] n13803_not ; n13804
g13549 and n13802_not n13803_not ; n13805
g13550 and n13804_not n13805_not ; n13806
g13551 and n13741_not n13752_not ; n13807
g13552 and n13738_not n13807_not ; n13808
g13553 and n13719_not n13725_not ; n13809
g13554 and b[55] n700 ; n13810
g13555 and b[53] n767 ; n13811
g13556 and b[54] n695 ; n13812
g13557 and n13811_not n13812_not ; n13813
g13558 and n13810_not n13813 ; n13814
g13559 and n703 n10684 ; n13815
g13560 and n13814 n13815_not ; n13816
g13561 and a[11] n13816_not ; n13817
g13562 and a[11] n13817_not ; n13818
g13563 and n13816_not n13817_not ; n13819
g13564 and n13818_not n13819_not ; n13820
g13565 and n13702_not n13705_not ; n13821
g13566 and b[52] n951 ; n13822
g13567 and b[50] n1056 ; n13823
g13568 and b[51] n946 ; n13824
g13569 and n13823_not n13824_not ; n13825
g13570 and n13822_not n13825 ; n13826
g13571 and n954 n9628 ; n13827
g13572 and n13826 n13827_not ; n13828
g13573 and a[14] n13828_not ; n13829
g13574 and a[14] n13829_not ; n13830
g13575 and n13828_not n13829_not ; n13831
g13576 and n13830_not n13831_not ; n13832
g13577 and n13694_not n13698_not ; n13833
g13578 and b[49] n1302 ; n13834
g13579 and b[47] n1391 ; n13835
g13580 and b[48] n1297 ; n13836
g13581 and n13835_not n13836_not ; n13837
g13582 and n13834_not n13837 ; n13838
g13583 and n1305 n8625 ; n13839
g13584 and n13838 n13839_not ; n13840
g13585 and a[17] n13840_not ; n13841
g13586 and a[17] n13841_not ; n13842
g13587 and n13840_not n13841_not ; n13843
g13588 and n13842_not n13843_not ; n13844
g13589 and n13686_not n13690_not ; n13845
g13590 and b[46] n1627 ; n13846
g13591 and b[44] n1763 ; n13847
g13592 and b[45] n1622 ; n13848
g13593 and n13847_not n13848_not ; n13849
g13594 and n13846_not n13849 ; n13850
g13595 and n1630 n7677 ; n13851
g13596 and n13850 n13851_not ; n13852
g13597 and a[20] n13852_not ; n13853
g13598 and a[20] n13853_not ; n13854
g13599 and n13852_not n13853_not ; n13855
g13600 and n13854_not n13855_not ; n13856
g13601 and n13678_not n13682_not ; n13857
g13602 and b[34] n3638 ; n13858
g13603 and b[32] n3843 ; n13859
g13604 and b[33] n3633 ; n13860
g13605 and n13859_not n13860_not ; n13861
g13606 and n13858_not n13861 ; n13862
g13607 and n3641 n4466 ; n13863
g13608 and n13862 n13863_not ; n13864
g13609 and a[32] n13864_not ; n13865
g13610 and a[32] n13865_not ; n13866
g13611 and n13864_not n13865_not ; n13867
g13612 and n13866_not n13867_not ; n13868
g13613 and b[22] n6595 ; n13869
g13614 and b[20] n6902 ; n13870
g13615 and b[21] n6590 ; n13871
g13616 and n13870_not n13871_not ; n13872
g13617 and n13869_not n13872 ; n13873
g13618 and n2145 n6598 ; n13874
g13619 and n13873 n13874_not ; n13875
g13620 and a[44] n13875_not ; n13876
g13621 and a[44] n13876_not ; n13877
g13622 and n13875_not n13876_not ; n13878
g13623 and n13877_not n13878_not ; n13879
g13624 and b[16] n8362 ; n13880
g13625 and b[14] n8715 ; n13881
g13626 and b[15] n8357 ; n13882
g13627 and n13881_not n13882_not ; n13883
g13628 and n13880_not n13883 ; n13884
g13629 and n1237 n8365 ; n13885
g13630 and n13884 n13885_not ; n13886
g13631 and a[50] n13886_not ; n13887
g13632 and a[50] n13887_not ; n13888
g13633 and n13886_not n13887_not ; n13889
g13634 and n13888_not n13889_not ; n13890
g13635 and b[10] n10426 ; n13891
g13636 and b[8] n10796 ; n13892
g13637 and b[9] n10421 ; n13893
g13638 and n13892_not n13893_not ; n13894
g13639 and n13891_not n13894 ; n13895
g13640 and n738 n10429 ; n13896
g13641 and n13895 n13896_not ; n13897
g13642 and a[56] n13897_not ; n13898
g13643 and a[56] n13898_not ; n13899
g13644 and n13897_not n13898_not ; n13900
g13645 and n13899_not n13900_not ; n13901
g13646 and n13521_not n13523_not ; n13902
g13647 and a[63] n13488 ; n13903
g13648 and b[0] n13903 ; n13904
g13649 and b[1] n13488_not ; n13905
g13650 and n13904_not n13905_not ; n13906
g13651 and b[4] n12668 ; n13907
g13652 and b[2] n13047 ; n13908
g13653 and b[3] n12663 ; n13909
g13654 and n13908_not n13909_not ; n13910
g13655 and n13907_not n13910 ; n13911
g13656 and n346 n12671 ; n13912
g13657 and n13911 n13912_not ; n13913
g13658 and a[62] n13913_not ; n13914
g13659 and a[62] n13914_not ; n13915
g13660 and n13913_not n13914_not ; n13916
g13661 and n13915_not n13916_not ; n13917
g13662 and n13906_not n13917_not ; n13918
g13663 and n13906_not n13918_not ; n13919
g13664 and n13917_not n13918_not ; n13920
g13665 and n13919_not n13920_not ; n13921
g13666 and n13490_not n13505_not ; n13922
g13667 and n13921 n13922 ; n13923
g13668 and n13921_not n13922_not ; n13924
g13669 and n13923_not n13924_not ; n13925
g13670 and b[7] n11531 ; n13926
g13671 and b[5] n11896 ; n13927
g13672 and b[6] n11526 ; n13928
g13673 and n13927_not n13928_not ; n13929
g13674 and n13926_not n13929 ; n13930
g13675 and n484 n11534 ; n13931
g13676 and n13930 n13931_not ; n13932
g13677 and a[59] n13932_not ; n13933
g13678 and a[59] n13933_not ; n13934
g13679 and n13932_not n13933_not ; n13935
g13680 and n13934_not n13935_not ; n13936
g13681 and n13925_not n13936 ; n13937
g13682 and n13925 n13936_not ; n13938
g13683 and n13937_not n13938_not ; n13939
g13684 and n13902_not n13939 ; n13940
g13685 and n13902 n13939_not ; n13941
g13686 and n13940_not n13941_not ; n13942
g13687 and n13901_not n13942 ; n13943
g13688 and n13942 n13943_not ; n13944
g13689 and n13901_not n13943_not ; n13945
g13690 and n13944_not n13945_not ; n13946
g13691 and n13474_not n13529_not ; n13947
g13692 and n13526_not n13947_not ; n13948
g13693 and n13946 n13948 ; n13949
g13694 and n13946_not n13948_not ; n13950
g13695 and n13949_not n13950_not ; n13951
g13696 and b[13] n9339 ; n13952
g13697 and b[11] n9732 ; n13953
g13698 and b[12] n9334 ; n13954
g13699 and n13953_not n13954_not ; n13955
g13700 and n13952_not n13955 ; n13956
g13701 and n1008 n9342 ; n13957
g13702 and n13956 n13957_not ; n13958
g13703 and a[53] n13958_not ; n13959
g13704 and a[53] n13959_not ; n13960
g13705 and n13958_not n13959_not ; n13961
g13706 and n13960_not n13961_not ; n13962
g13707 and n13951_not n13962 ; n13963
g13708 and n13951 n13962_not ; n13964
g13709 and n13963_not n13964_not ; n13965
g13710 and n13545_not n13547_not ; n13966
g13711 and n13965 n13966_not ; n13967
g13712 and n13965_not n13966 ; n13968
g13713 and n13967_not n13968_not ; n13969
g13714 and n13890_not n13969 ; n13970
g13715 and n13969 n13970_not ; n13971
g13716 and n13890_not n13970_not ; n13972
g13717 and n13971_not n13972_not ; n13973
g13718 and n13550_not n13556_not ; n13974
g13719 and n13973 n13974 ; n13975
g13720 and n13973_not n13974_not ; n13976
g13721 and n13975_not n13976_not ; n13977
g13722 and b[19] n7446 ; n13978
g13723 and b[17] n7787 ; n13979
g13724 and b[18] n7441 ; n13980
g13725 and n13979_not n13980_not ; n13981
g13726 and n13978_not n13981 ; n13982
g13727 and n1708 n7449 ; n13983
g13728 and n13982 n13983_not ; n13984
g13729 and a[47] n13984_not ; n13985
g13730 and a[47] n13985_not ; n13986
g13731 and n13984_not n13985_not ; n13987
g13732 and n13986_not n13987_not ; n13988
g13733 and n13977_not n13988 ; n13989
g13734 and n13977 n13988_not ; n13990
g13735 and n13989_not n13990_not ; n13991
g13736 and n13570_not n13572_not ; n13992
g13737 and n13991 n13992_not ; n13993
g13738 and n13991_not n13992 ; n13994
g13739 and n13993_not n13994_not ; n13995
g13740 and n13879_not n13995 ; n13996
g13741 and n13995 n13996_not ; n13997
g13742 and n13879_not n13996_not ; n13998
g13743 and n13997_not n13998_not ; n13999
g13744 and n13575_not n13578_not ; n14000
g13745 and n13999 n14000 ; n14001
g13746 and n13999_not n14000_not ; n14002
g13747 and n14001_not n14002_not ; n14003
g13748 and b[25] n5777 ; n14004
g13749 and b[23] n6059 ; n14005
g13750 and b[24] n5772 ; n14006
g13751 and n14005_not n14006_not ; n14007
g13752 and n14004_not n14007 ; n14008
g13753 and n2485 n5780 ; n14009
g13754 and n14008 n14009_not ; n14010
g13755 and a[41] n14010_not ; n14011
g13756 and a[41] n14011_not ; n14012
g13757 and n14010_not n14011_not ; n14013
g13758 and n14012_not n14013_not ; n14014
g13759 and n14003 n14014_not ; n14015
g13760 and n14003 n14015_not ; n14016
g13761 and n14014_not n14015_not ; n14017
g13762 and n14016_not n14017_not ; n14018
g13763 and n13592_not n13598_not ; n14019
g13764 and n14018 n14019 ; n14020
g13765 and n14018_not n14019_not ; n14021
g13766 and n14020_not n14021_not ; n14022
g13767 and b[28] n5035 ; n14023
g13768 and b[26] n5277 ; n14024
g13769 and b[27] n5030 ; n14025
g13770 and n14024_not n14025_not ; n14026
g13771 and n14023_not n14026 ; n14027
g13772 and n3189 n5038 ; n14028
g13773 and n14027 n14028_not ; n14029
g13774 and a[38] n14029_not ; n14030
g13775 and a[38] n14030_not ; n14031
g13776 and n14029_not n14030_not ; n14032
g13777 and n14031_not n14032_not ; n14033
g13778 and n14022 n14033_not ; n14034
g13779 and n14022 n14034_not ; n14035
g13780 and n14033_not n14034_not ; n14036
g13781 and n14035_not n14036_not ; n14037
g13782 and n13611_not n13617_not ; n14038
g13783 and n14037 n14038 ; n14039
g13784 and n14037_not n14038_not ; n14040
g13785 and n14039_not n14040_not ; n14041
g13786 and b[31] n4287 ; n14042
g13787 and b[29] n4532 ; n14043
g13788 and b[30] n4282 ; n14044
g13789 and n14043_not n14044_not ; n14045
g13790 and n14042_not n14045 ; n14046
g13791 and n3796 n4290 ; n14047
g13792 and n14046 n14047_not ; n14048
g13793 and a[35] n14048_not ; n14049
g13794 and a[35] n14049_not ; n14050
g13795 and n14048_not n14049_not ; n14051
g13796 and n14050_not n14051_not ; n14052
g13797 and n14041_not n14052 ; n14053
g13798 and n14041 n14052_not ; n14054
g13799 and n14053_not n14054_not ; n14055
g13800 and n13631_not n13634_not ; n14056
g13801 and n14055 n14056_not ; n14057
g13802 and n14055_not n14056 ; n14058
g13803 and n14057_not n14058_not ; n14059
g13804 and n13868_not n14059 ; n14060
g13805 and n14059 n14060_not ; n14061
g13806 and n13868_not n14060_not ; n14062
g13807 and n14061_not n14062_not ; n14063
g13808 and n13207_not n13640_not ; n14064
g13809 and n13637_not n14064_not ; n14065
g13810 and n14063 n14065 ; n14066
g13811 and n14063_not n14065_not ; n14067
g13812 and n14066_not n14067_not ; n14068
g13813 and b[37] n3050 ; n14069
g13814 and b[35] n3243 ; n14070
g13815 and b[36] n3045 ; n14071
g13816 and n14070_not n14071_not ; n14072
g13817 and n14069_not n14072 ; n14073
g13818 and n3053 n5181 ; n14074
g13819 and n14073 n14074_not ; n14075
g13820 and a[29] n14075_not ; n14076
g13821 and a[29] n14076_not ; n14077
g13822 and n14075_not n14076_not ; n14078
g13823 and n14077_not n14078_not ; n14079
g13824 and n14068 n14079_not ; n14080
g13825 and n14068 n14080_not ; n14081
g13826 and n14079_not n14080_not ; n14082
g13827 and n14081_not n14082_not ; n14083
g13828 and n13655_not n13659_not ; n14084
g13829 and n14083 n14084 ; n14085
g13830 and n14083_not n14084_not ; n14086
g13831 and n14085_not n14086_not ; n14087
g13832 and b[40] n2539 ; n14088
g13833 and b[38] n2685 ; n14089
g13834 and b[39] n2534 ; n14090
g13835 and n14089_not n14090_not ; n14091
g13836 and n14088_not n14091 ; n14092
g13837 and n2542 n5955 ; n14093
g13838 and n14092 n14093_not ; n14094
g13839 and a[26] n14094_not ; n14095
g13840 and a[26] n14095_not ; n14096
g13841 and n14094_not n14095_not ; n14097
g13842 and n14096_not n14097_not ; n14098
g13843 and n14087 n14098_not ; n14099
g13844 and n14087 n14099_not ; n14100
g13845 and n14098_not n14099_not ; n14101
g13846 and n14100_not n14101_not ; n14102
g13847 and n13673_not n13675_not ; n14103
g13848 and n14102_not n14103_not ; n14104
g13849 and n14102_not n14104_not ; n14105
g13850 and n14103_not n14104_not ; n14106
g13851 and n14105_not n14106_not ; n14107
g13852 and b[43] n2048 ; n14108
g13853 and b[41] n2198 ; n14109
g13854 and b[42] n2043 ; n14110
g13855 and n14109_not n14110_not ; n14111
g13856 and n14108_not n14111 ; n14112
g13857 and n2051 n6515 ; n14113
g13858 and n14112 n14113_not ; n14114
g13859 and a[23] n14114_not ; n14115
g13860 and a[23] n14115_not ; n14116
g13861 and n14114_not n14115_not ; n14117
g13862 and n14116_not n14117_not ; n14118
g13863 and n14107_not n14118 ; n14119
g13864 and n14107 n14118_not ; n14120
g13865 and n14119_not n14120_not ; n14121
g13866 and n13857_not n14121_not ; n14122
g13867 and n13857 n14121 ; n14123
g13868 and n14122_not n14123_not ; n14124
g13869 and n13856_not n14124 ; n14125
g13870 and n13856_not n14125_not ; n14126
g13871 and n14124 n14125_not ; n14127
g13872 and n14126_not n14127_not ; n14128
g13873 and n13845_not n14128_not ; n14129
g13874 and n13845 n14127_not ; n14130
g13875 and n14126_not n14130 ; n14131
g13876 and n14129_not n14131_not ; n14132
g13877 and n13844_not n14132 ; n14133
g13878 and n13844_not n14133_not ; n14134
g13879 and n14132 n14133_not ; n14135
g13880 and n14134_not n14135_not ; n14136
g13881 and n13833_not n14136_not ; n14137
g13882 and n13833 n14135_not ; n14138
g13883 and n14134_not n14138 ; n14139
g13884 and n14137_not n14139_not ; n14140
g13885 and n13832_not n14140 ; n14141
g13886 and n13832 n14140_not ; n14142
g13887 and n14141_not n14142_not ; n14143
g13888 and n13821_not n14143 ; n14144
g13889 and n13821 n14143_not ; n14145
g13890 and n14144_not n14145_not ; n14146
g13891 and n13820_not n14146 ; n14147
g13892 and n13820 n14146_not ; n14148
g13893 and n14147_not n14148_not ; n14149
g13894 and n13809_not n14149 ; n14150
g13895 and n13809 n14149_not ; n14151
g13896 and n14150_not n14151_not ; n14152
g13897 and b[58] n511 ; n14153
g13898 and b[56] n541 ; n14154
g13899 and b[57] n506 ; n14155
g13900 and n14154_not n14155_not ; n14156
g13901 and n14153_not n14156 ; n14157
g13902 and n514 n11436 ; n14158
g13903 and n14157 n14158_not ; n14159
g13904 and a[8] n14159_not ; n14160
g13905 and a[8] n14160_not ; n14161
g13906 and n14159_not n14160_not ; n14162
g13907 and n14161_not n14162_not ; n14163
g13908 and n14152 n14163_not ; n14164
g13909 and n14152 n14164_not ; n14165
g13910 and n14163_not n14164_not ; n14166
g13911 and n14165_not n14166_not ; n14167
g13912 and b[61] n362 ; n14168
g13913 and b[59] n403 ; n14169
g13914 and b[60] n357 ; n14170
g13915 and n14169_not n14170_not ; n14171
g13916 and n14168_not n14171 ; n14172
g13917 and n365 n12969 ; n14173
g13918 and n14172 n14173_not ; n14174
g13919 and a[5] n14174_not ; n14175
g13920 and a[5] n14175_not ; n14176
g13921 and n14174_not n14175_not ; n14177
g13922 and n14176_not n14177_not ; n14178
g13923 and n14167_not n14178 ; n14179
g13924 and n14167 n14178_not ; n14180
g13925 and n14179_not n14180_not ; n14181
g13926 and n13808_not n14181_not ; n14182
g13927 and n13808 n14181 ; n14183
g13928 and n14182_not n14183_not ; n14184
g13929 and n13806_not n14184 ; n14185
g13930 and n13806 n14184_not ; n14186
g13931 and n14185_not n14186_not ; n14187
g13932 and n13792_not n14187 ; n14188
g13933 and n13792 n14187_not ; n14189
g13934 and n14188_not n14189_not ; n14190
g13935 and n13791_not n14190 ; n14191
g13936 and n13791 n14190_not ; n14192
g13937 and n14191_not n14192_not ; f[64]
g13938 and b[53] n951 ; n14194
g13939 and b[51] n1056 ; n14195
g13940 and b[52] n946 ; n14196
g13941 and n14195_not n14196_not ; n14197
g13942 and n14194_not n14197 ; n14198
g13943 and n954 n9972 ; n14199
g13944 and n14198 n14199_not ; n14200
g13945 and a[14] n14200_not ; n14201
g13946 and a[14] n14201_not ; n14202
g13947 and n14200_not n14201_not ; n14203
g13948 and n14202_not n14203_not ; n14204
g13949 and n14133_not n14137_not ; n14205
g13950 and n14125_not n14129_not ; n14206
g13951 and b[47] n1627 ; n14207
g13952 and b[45] n1763 ; n14208
g13953 and b[46] n1622 ; n14209
g13954 and n14208_not n14209_not ; n14210
g13955 and n14207_not n14210 ; n14211
g13956 and n1630 n7703 ; n14212
g13957 and n14211 n14212_not ; n14213
g13958 and a[20] n14213_not ; n14214
g13959 and a[20] n14214_not ; n14215
g13960 and n14213_not n14214_not ; n14216
g13961 and n14215_not n14216_not ; n14217
g13962 and n14099_not n14104_not ; n14218
g13963 and n14054_not n14057_not ; n14219
g13964 and n13996_not n14002_not ; n14220
g13965 and n13990_not n13993_not ; n14221
g13966 and n13970_not n13976_not ; n14222
g13967 and n13964_not n13967_not ; n14223
g13968 and b[14] n9339 ; n14224
g13969 and b[12] n9732 ; n14225
g13970 and b[13] n9334 ; n14226
g13971 and n14225_not n14226_not ; n14227
g13972 and n14224_not n14227 ; n14228
g13973 and n1034 n9342 ; n14229
g13974 and n14228 n14229_not ; n14230
g13975 and a[53] n14230_not ; n14231
g13976 and a[53] n14231_not ; n14232
g13977 and n14230_not n14231_not ; n14233
g13978 and n14232_not n14233_not ; n14234
g13979 and n13943_not n13950_not ; n14235
g13980 and n13938_not n13940_not ; n14236
g13981 and b[1] n13903 ; n14237
g13982 and b[2] n13488_not ; n14238
g13983 and n14237_not n14238_not ; n14239
g13984 and b[5] n12668 ; n14240
g13985 and b[3] n13047 ; n14241
g13986 and b[4] n12663 ; n14242
g13987 and n14241_not n14242_not ; n14243
g13988 and n14240_not n14243 ; n14244
g13989 and n394 n12671 ; n14245
g13990 and n14244 n14245_not ; n14246
g13991 and a[62] n14246_not ; n14247
g13992 and a[62] n14247_not ; n14248
g13993 and n14246_not n14247_not ; n14249
g13994 and n14248_not n14249_not ; n14250
g13995 and n14239_not n14250_not ; n14251
g13996 and n14239_not n14251_not ; n14252
g13997 and n14250_not n14251_not ; n14253
g13998 and n14252_not n14253_not ; n14254
g13999 and n13918_not n13924_not ; n14255
g14000 and n14254 n14255 ; n14256
g14001 and n14254_not n14255_not ; n14257
g14002 and n14256_not n14257_not ; n14258
g14003 and b[8] n11531 ; n14259
g14004 and b[6] n11896 ; n14260
g14005 and b[7] n11526 ; n14261
g14006 and n14260_not n14261_not ; n14262
g14007 and n14259_not n14262 ; n14263
g14008 and n585 n11534 ; n14264
g14009 and n14263 n14264_not ; n14265
g14010 and a[59] n14265_not ; n14266
g14011 and a[59] n14266_not ; n14267
g14012 and n14265_not n14266_not ; n14268
g14013 and n14267_not n14268_not ; n14269
g14014 and n14258 n14269_not ; n14270
g14015 and n14258_not n14269 ; n14271
g14016 and n14236_not n14271_not ; n14272
g14017 and n14270_not n14272 ; n14273
g14018 and n14236_not n14273_not ; n14274
g14019 and n14270_not n14273_not ; n14275
g14020 and n14271_not n14275 ; n14276
g14021 and n14274_not n14276_not ; n14277
g14022 and b[11] n10426 ; n14278
g14023 and b[9] n10796 ; n14279
g14024 and b[10] n10421 ; n14280
g14025 and n14279_not n14280_not ; n14281
g14026 and n14278_not n14281 ; n14282
g14027 and n818 n10429 ; n14283
g14028 and n14282 n14283_not ; n14284
g14029 and a[56] n14284_not ; n14285
g14030 and a[56] n14285_not ; n14286
g14031 and n14284_not n14285_not ; n14287
g14032 and n14286_not n14287_not ; n14288
g14033 and n14277 n14288 ; n14289
g14034 and n14277_not n14288_not ; n14290
g14035 and n14289_not n14290_not ; n14291
g14036 and n14235_not n14291 ; n14292
g14037 and n14235 n14291_not ; n14293
g14038 and n14292_not n14293_not ; n14294
g14039 and n14234_not n14294 ; n14295
g14040 and n14294 n14295_not ; n14296
g14041 and n14234_not n14295_not ; n14297
g14042 and n14296_not n14297_not ; n14298
g14043 and n14223_not n14298 ; n14299
g14044 and n14223 n14298_not ; n14300
g14045 and n14299_not n14300_not ; n14301
g14046 and b[17] n8362 ; n14302
g14047 and b[15] n8715 ; n14303
g14048 and b[16] n8357 ; n14304
g14049 and n14303_not n14304_not ; n14305
g14050 and n14302_not n14305 ; n14306
g14051 and n1356 n8365 ; n14307
g14052 and n14306 n14307_not ; n14308
g14053 and a[50] n14308_not ; n14309
g14054 and a[50] n14309_not ; n14310
g14055 and n14308_not n14309_not ; n14311
g14056 and n14310_not n14311_not ; n14312
g14057 and n14301_not n14312_not ; n14313
g14058 and n14301 n14312 ; n14314
g14059 and n14313_not n14314_not ; n14315
g14060 and n14222 n14315_not ; n14316
g14061 and n14222_not n14315 ; n14317
g14062 and n14316_not n14317_not ; n14318
g14063 and b[20] n7446 ; n14319
g14064 and b[18] n7787 ; n14320
g14065 and b[19] n7441 ; n14321
g14066 and n14320_not n14321_not ; n14322
g14067 and n14319_not n14322 ; n14323
g14068 and n1846 n7449 ; n14324
g14069 and n14323 n14324_not ; n14325
g14070 and a[47] n14325_not ; n14326
g14071 and a[47] n14326_not ; n14327
g14072 and n14325_not n14326_not ; n14328
g14073 and n14327_not n14328_not ; n14329
g14074 and n14318 n14329_not ; n14330
g14075 and n14318 n14330_not ; n14331
g14076 and n14329_not n14330_not ; n14332
g14077 and n14331_not n14332_not ; n14333
g14078 and n14221_not n14333 ; n14334
g14079 and n14221 n14333_not ; n14335
g14080 and n14334_not n14335_not ; n14336
g14081 and b[23] n6595 ; n14337
g14082 and b[21] n6902 ; n14338
g14083 and b[22] n6590 ; n14339
g14084 and n14338_not n14339_not ; n14340
g14085 and n14337_not n14340 ; n14341
g14086 and n2300 n6598 ; n14342
g14087 and n14341 n14342_not ; n14343
g14088 and a[44] n14343_not ; n14344
g14089 and a[44] n14344_not ; n14345
g14090 and n14343_not n14344_not ; n14346
g14091 and n14345_not n14346_not ; n14347
g14092 and n14336_not n14347_not ; n14348
g14093 and n14336 n14347 ; n14349
g14094 and n14348_not n14349_not ; n14350
g14095 and n14220 n14350_not ; n14351
g14096 and n14220_not n14350 ; n14352
g14097 and n14351_not n14352_not ; n14353
g14098 and b[26] n5777 ; n14354
g14099 and b[24] n6059 ; n14355
g14100 and b[25] n5772 ; n14356
g14101 and n14355_not n14356_not ; n14357
g14102 and n14354_not n14357 ; n14358
g14103 and n2813 n5780 ; n14359
g14104 and n14358 n14359_not ; n14360
g14105 and a[41] n14360_not ; n14361
g14106 and a[41] n14361_not ; n14362
g14107 and n14360_not n14361_not ; n14363
g14108 and n14362_not n14363_not ; n14364
g14109 and n14353 n14364_not ; n14365
g14110 and n14353 n14365_not ; n14366
g14111 and n14364_not n14365_not ; n14367
g14112 and n14366_not n14367_not ; n14368
g14113 and n14015_not n14021_not ; n14369
g14114 and n14368 n14369 ; n14370
g14115 and n14368_not n14369_not ; n14371
g14116 and n14370_not n14371_not ; n14372
g14117 and b[29] n5035 ; n14373
g14118 and b[27] n5277 ; n14374
g14119 and b[28] n5030 ; n14375
g14120 and n14374_not n14375_not ; n14376
g14121 and n14373_not n14376 ; n14377
g14122 and n3383 n5038 ; n14378
g14123 and n14377 n14378_not ; n14379
g14124 and a[38] n14379_not ; n14380
g14125 and a[38] n14380_not ; n14381
g14126 and n14379_not n14380_not ; n14382
g14127 and n14381_not n14382_not ; n14383
g14128 and n14372 n14383_not ; n14384
g14129 and n14372 n14384_not ; n14385
g14130 and n14383_not n14384_not ; n14386
g14131 and n14385_not n14386_not ; n14387
g14132 and n14034_not n14040_not ; n14388
g14133 and n14387 n14388 ; n14389
g14134 and n14387_not n14388_not ; n14390
g14135 and n14389_not n14390_not ; n14391
g14136 and b[32] n4287 ; n14392
g14137 and b[30] n4532 ; n14393
g14138 and b[31] n4282 ; n14394
g14139 and n14393_not n14394_not ; n14395
g14140 and n14392_not n14395 ; n14396
g14141 and n4013 n4290 ; n14397
g14142 and n14396 n14397_not ; n14398
g14143 and a[35] n14398_not ; n14399
g14144 and a[35] n14399_not ; n14400
g14145 and n14398_not n14399_not ; n14401
g14146 and n14400_not n14401_not ; n14402
g14147 and n14391 n14402_not ; n14403
g14148 and n14391_not n14402 ; n14404
g14149 and n14219_not n14404_not ; n14405
g14150 and n14403_not n14405 ; n14406
g14151 and n14219_not n14406_not ; n14407
g14152 and n14403_not n14406_not ; n14408
g14153 and n14404_not n14408 ; n14409
g14154 and n14407_not n14409_not ; n14410
g14155 and b[35] n3638 ; n14411
g14156 and b[33] n3843 ; n14412
g14157 and b[34] n3633 ; n14413
g14158 and n14412_not n14413_not ; n14414
g14159 and n14411_not n14414 ; n14415
g14160 and n3641 n4696 ; n14416
g14161 and n14415 n14416_not ; n14417
g14162 and a[32] n14417_not ; n14418
g14163 and a[32] n14418_not ; n14419
g14164 and n14417_not n14418_not ; n14420
g14165 and n14419_not n14420_not ; n14421
g14166 and n14410_not n14421_not ; n14422
g14167 and n14410_not n14422_not ; n14423
g14168 and n14421_not n14422_not ; n14424
g14169 and n14423_not n14424_not ; n14425
g14170 and n14060_not n14067_not ; n14426
g14171 and n14425 n14426 ; n14427
g14172 and n14425_not n14426_not ; n14428
g14173 and n14427_not n14428_not ; n14429
g14174 and b[38] n3050 ; n14430
g14175 and b[36] n3243 ; n14431
g14176 and b[37] n3045 ; n14432
g14177 and n14431_not n14432_not ; n14433
g14178 and n14430_not n14433 ; n14434
g14179 and n3053 n5205 ; n14435
g14180 and n14434 n14435_not ; n14436
g14181 and a[29] n14436_not ; n14437
g14182 and a[29] n14437_not ; n14438
g14183 and n14436_not n14437_not ; n14439
g14184 and n14438_not n14439_not ; n14440
g14185 and n14429 n14440_not ; n14441
g14186 and n14429 n14441_not ; n14442
g14187 and n14440_not n14441_not ; n14443
g14188 and n14442_not n14443_not ; n14444
g14189 and n14080_not n14086_not ; n14445
g14190 and n14444 n14445 ; n14446
g14191 and n14444_not n14445_not ; n14447
g14192 and n14446_not n14447_not ; n14448
g14193 and b[41] n2539 ; n14449
g14194 and b[39] n2685 ; n14450
g14195 and b[40] n2534 ; n14451
g14196 and n14450_not n14451_not ; n14452
g14197 and n14449_not n14452 ; n14453
g14198 and n2542 n6219 ; n14454
g14199 and n14453 n14454_not ; n14455
g14200 and a[26] n14455_not ; n14456
g14201 and a[26] n14456_not ; n14457
g14202 and n14455_not n14456_not ; n14458
g14203 and n14457_not n14458_not ; n14459
g14204 and n14448 n14459_not ; n14460
g14205 and n14448_not n14459 ; n14461
g14206 and n14218_not n14461_not ; n14462
g14207 and n14460_not n14462 ; n14463
g14208 and n14218_not n14463_not ; n14464
g14209 and n14460_not n14463_not ; n14465
g14210 and n14461_not n14465 ; n14466
g14211 and n14464_not n14466_not ; n14467
g14212 and b[44] n2048 ; n14468
g14213 and b[42] n2198 ; n14469
g14214 and b[43] n2043 ; n14470
g14215 and n14469_not n14470_not ; n14471
g14216 and n14468_not n14471 ; n14472
g14217 and n2051 n7072 ; n14473
g14218 and n14472 n14473_not ; n14474
g14219 and a[23] n14474_not ; n14475
g14220 and a[23] n14475_not ; n14476
g14221 and n14474_not n14475_not ; n14477
g14222 and n14476_not n14477_not ; n14478
g14223 and n14467_not n14478_not ; n14479
g14224 and n14467_not n14479_not ; n14480
g14225 and n14478_not n14479_not ; n14481
g14226 and n14480_not n14481_not ; n14482
g14227 and n14107_not n14118_not ; n14483
g14228 and n14122_not n14483_not ; n14484
g14229 and n14482_not n14484_not ; n14485
g14230 and n14482 n14484 ; n14486
g14231 and n14485_not n14486_not ; n14487
g14232 and n14217_not n14487 ; n14488
g14233 and n14217_not n14488_not ; n14489
g14234 and n14487 n14488_not ; n14490
g14235 and n14489_not n14490_not ; n14491
g14236 and n14206_not n14491_not ; n14492
g14237 and n14206_not n14492_not ; n14493
g14238 and n14491_not n14492_not ; n14494
g14239 and n14493_not n14494_not ; n14495
g14240 and b[50] n1302 ; n14496
g14241 and b[48] n1391 ; n14497
g14242 and b[49] n1297 ; n14498
g14243 and n14497_not n14498_not ; n14499
g14244 and n14496_not n14499 ; n14500
g14245 and n1305 n8949 ; n14501
g14246 and n14500 n14501_not ; n14502
g14247 and a[17] n14502_not ; n14503
g14248 and a[17] n14503_not ; n14504
g14249 and n14502_not n14503_not ; n14505
g14250 and n14504_not n14505_not ; n14506
g14251 and n14495 n14506 ; n14507
g14252 and n14495_not n14506_not ; n14508
g14253 and n14507_not n14508_not ; n14509
g14254 and n14205_not n14509 ; n14510
g14255 and n14205 n14509_not ; n14511
g14256 and n14510_not n14511_not ; n14512
g14257 and n14204_not n14512 ; n14513
g14258 and n14512 n14513_not ; n14514
g14259 and n14204_not n14513_not ; n14515
g14260 and n14514_not n14515_not ; n14516
g14261 and n14141_not n14144_not ; n14517
g14262 and n14516 n14517 ; n14518
g14263 and n14516_not n14517_not ; n14519
g14264 and n14518_not n14519_not ; n14520
g14265 and b[56] n700 ; n14521
g14266 and b[54] n767 ; n14522
g14267 and b[55] n695 ; n14523
g14268 and n14522_not n14523_not ; n14524
g14269 and n14521_not n14524 ; n14525
g14270 and n703 n10708 ; n14526
g14271 and n14525 n14526_not ; n14527
g14272 and a[11] n14527_not ; n14528
g14273 and a[11] n14528_not ; n14529
g14274 and n14527_not n14528_not ; n14530
g14275 and n14529_not n14530_not ; n14531
g14276 and n14520_not n14531 ; n14532
g14277 and n14520 n14531_not ; n14533
g14278 and n14532_not n14533_not ; n14534
g14279 and b[59] n511 ; n14535
g14280 and b[57] n541 ; n14536
g14281 and b[58] n506 ; n14537
g14282 and n14536_not n14537_not ; n14538
g14283 and n14535_not n14538 ; n14539
g14284 and n514 n12179 ; n14540
g14285 and n14539 n14540_not ; n14541
g14286 and a[8] n14541_not ; n14542
g14287 and a[8] n14542_not ; n14543
g14288 and n14541_not n14542_not ; n14544
g14289 and n14543_not n14544_not ; n14545
g14290 and n14534 n14545_not ; n14546
g14291 and n14534 n14546_not ; n14547
g14292 and n14545_not n14546_not ; n14548
g14293 and n14547_not n14548_not ; n14549
g14294 and n14147_not n14150_not ; n14550
g14295 and n14549 n14550 ; n14551
g14296 and n14549_not n14550_not ; n14552
g14297 and n14551_not n14552_not ; n14553
g14298 and b[62] n362 ; n14554
g14299 and b[60] n403 ; n14555
g14300 and b[61] n357 ; n14556
g14301 and n14555_not n14556_not ; n14557
g14302 and n14554_not n14557 ; n14558
g14303 and n365 n13370 ; n14559
g14304 and n14558 n14559_not ; n14560
g14305 and a[5] n14560_not ; n14561
g14306 and a[5] n14561_not ; n14562
g14307 and n14560_not n14561_not ; n14563
g14308 and n14562_not n14563_not ; n14564
g14309 and n14553 n14564_not ; n14565
g14310 and n14553 n14565_not ; n14566
g14311 and n14564_not n14565_not ; n14567
g14312 and n14566_not n14567_not ; n14568
g14313 and n14167_not n14178_not ; n14569
g14314 and n14164_not n14569_not ; n14570
g14315 and n269 n13797 ; n14571
g14316 and a[2]_not n14571_not ; n14572
g14317 and b[63] n284 ; n14573
g14318 and n14571_not n14573_not ; n14574
g14319 and a[2] n14574_not ; n14575
g14320 and n14572_not n14575_not ; n14576
g14321 and n14570_not n14576 ; n14577
g14322 and n14570 n14576_not ; n14578
g14323 and n14577_not n14578_not ; n14579
g14324 and n14568_not n14579 ; n14580
g14325 and n14568_not n14580_not ; n14581
g14326 and n14579 n14580_not ; n14582
g14327 and n14581_not n14582_not ; n14583
g14328 and n14182_not n14185_not ; n14584
g14329 and n14583 n14584 ; n14585
g14330 and n14583_not n14584_not ; n14586
g14331 and n14585_not n14586_not ; n14587
g14332 and n14188_not n14191_not ; n14588
g14333 and n14587 n14588_not ; n14589
g14334 and n14587_not n14588 ; n14590
g14335 and n14589_not n14590_not ; f[65]
g14336 and n14552_not n14565_not ; n14592
g14337 and b[63] n362 ; n14593
g14338 and b[61] n403 ; n14594
g14339 and b[62] n357 ; n14595
g14340 and n14594_not n14595_not ; n14596
g14341 and n14593_not n14596 ; n14597
g14342 and n365 n13771 ; n14598
g14343 and n14597 n14598_not ; n14599
g14344 and a[5] n14599_not ; n14600
g14345 and a[5] n14600_not ; n14601
g14346 and n14599_not n14600_not ; n14602
g14347 and n14601_not n14602_not ; n14603
g14348 and n14592_not n14603_not ; n14604
g14349 and n14592_not n14604_not ; n14605
g14350 and n14603_not n14604_not ; n14606
g14351 and n14605_not n14606_not ; n14607
g14352 and b[57] n700 ; n14608
g14353 and b[55] n767 ; n14609
g14354 and b[56] n695 ; n14610
g14355 and n14609_not n14610_not ; n14611
g14356 and n14608_not n14611 ; n14612
g14357 and n703 n11410 ; n14613
g14358 and n14612 n14613_not ; n14614
g14359 and a[11] n14614_not ; n14615
g14360 and a[11] n14615_not ; n14616
g14361 and n14614_not n14615_not ; n14617
g14362 and n14616_not n14617_not ; n14618
g14363 and n14513_not n14519_not ; n14619
g14364 and n14618 n14619 ; n14620
g14365 and n14618_not n14619_not ; n14621
g14366 and n14620_not n14621_not ; n14622
g14367 and b[51] n1302 ; n14623
g14368 and b[49] n1391 ; n14624
g14369 and b[50] n1297 ; n14625
g14370 and n14624_not n14625_not ; n14626
g14371 and n14623_not n14626 ; n14627
g14372 and n1305 n8976 ; n14628
g14373 and n14627 n14628_not ; n14629
g14374 and a[17] n14629_not ; n14630
g14375 and a[17] n14630_not ; n14631
g14376 and n14629_not n14630_not ; n14632
g14377 and n14631_not n14632_not ; n14633
g14378 and n14488_not n14492_not ; n14634
g14379 and n14633 n14634 ; n14635
g14380 and n14633_not n14634_not ; n14636
g14381 and n14635_not n14636_not ; n14637
g14382 and b[48] n1627 ; n14638
g14383 and b[46] n1763 ; n14639
g14384 and b[47] n1622 ; n14640
g14385 and n14639_not n14640_not ; n14641
g14386 and n14638_not n14641 ; n14642
g14387 and n1630 n8009 ; n14643
g14388 and n14642 n14643_not ; n14644
g14389 and a[20] n14644_not ; n14645
g14390 and a[20] n14645_not ; n14646
g14391 and n14644_not n14645_not ; n14647
g14392 and n14646_not n14647_not ; n14648
g14393 and n14479_not n14485_not ; n14649
g14394 and n14648 n14649 ; n14650
g14395 and n14648_not n14649_not ; n14651
g14396 and n14650_not n14651_not ; n14652
g14397 and b[45] n2048 ; n14653
g14398 and b[43] n2198 ; n14654
g14399 and b[44] n2043 ; n14655
g14400 and n14654_not n14655_not ; n14656
g14401 and n14653_not n14656 ; n14657
g14402 and n2051 n7361 ; n14658
g14403 and n14657 n14658_not ; n14659
g14404 and a[23] n14659_not ; n14660
g14405 and a[23] n14660_not ; n14661
g14406 and n14659_not n14660_not ; n14662
g14407 and n14661_not n14662_not ; n14663
g14408 and n14465_not n14663 ; n14664
g14409 and n14465 n14663_not ; n14665
g14410 and n14664_not n14665_not ; n14666
g14411 and b[42] n2539 ; n14667
g14412 and b[40] n2685 ; n14668
g14413 and b[41] n2534 ; n14669
g14414 and n14668_not n14669_not ; n14670
g14415 and n14667_not n14670 ; n14671
g14416 and n2542 n6489 ; n14672
g14417 and n14671 n14672_not ; n14673
g14418 and a[26] n14673_not ; n14674
g14419 and a[26] n14674_not ; n14675
g14420 and n14673_not n14674_not ; n14676
g14421 and n14675_not n14676_not ; n14677
g14422 and n14441_not n14447_not ; n14678
g14423 and n14677 n14678 ; n14679
g14424 and n14677_not n14678_not ; n14680
g14425 and n14679_not n14680_not ; n14681
g14426 and n14422_not n14428_not ; n14682
g14427 and b[39] n3050 ; n14683
g14428 and b[37] n3243 ; n14684
g14429 and b[38] n3045 ; n14685
g14430 and n14684_not n14685_not ; n14686
g14431 and n14683_not n14686 ; n14687
g14432 and n3053_not n14687 ; n14688
g14433 and n5451_not n14687 ; n14689
g14434 and n14688_not n14689_not ; n14690
g14435 and a[29] n14690_not ; n14691
g14436 and a[29]_not n14690 ; n14692
g14437 and n14691_not n14692_not ; n14693
g14438 and n14682_not n14693_not ; n14694
g14439 and n14682 n14693 ; n14695
g14440 and n14694_not n14695_not ; n14696
g14441 and b[33] n4287 ; n14697
g14442 and b[31] n4532 ; n14698
g14443 and b[32] n4282 ; n14699
g14444 and n14698_not n14699_not ; n14700
g14445 and n14697_not n14700 ; n14701
g14446 and n4223 n4290 ; n14702
g14447 and n14701 n14702_not ; n14703
g14448 and a[35] n14703_not ; n14704
g14449 and a[35] n14704_not ; n14705
g14450 and n14703_not n14704_not ; n14706
g14451 and n14705_not n14706_not ; n14707
g14452 and b[24] n6595 ; n14708
g14453 and b[22] n6902 ; n14709
g14454 and b[23] n6590 ; n14710
g14455 and n14709_not n14710_not ; n14711
g14456 and n14708_not n14711 ; n14712
g14457 and n2458 n6598 ; n14713
g14458 and n14712 n14713_not ; n14714
g14459 and a[44] n14714_not ; n14715
g14460 and a[44] n14715_not ; n14716
g14461 and n14714_not n14715_not ; n14717
g14462 and n14716_not n14717_not ; n14718
g14463 and b[15] n9339 ; n14719
g14464 and b[13] n9732 ; n14720
g14465 and b[14] n9334 ; n14721
g14466 and n14720_not n14721_not ; n14722
g14467 and n14719_not n14722 ; n14723
g14468 and n1131 n9342 ; n14724
g14469 and n14723 n14724_not ; n14725
g14470 and a[53] n14725_not ; n14726
g14471 and a[53] n14726_not ; n14727
g14472 and n14725_not n14726_not ; n14728
g14473 and n14727_not n14728_not ; n14729
g14474 and n14290_not n14292_not ; n14730
g14475 and n14251_not n14257_not ; n14731
g14476 and b[2] n13903 ; n14732
g14477 and b[3] n13488_not ; n14733
g14478 and n14732_not n14733_not ; n14734
g14479 and a[2] n14734_not ; n14735
g14480 and a[2]_not n14734 ; n14736
g14481 and n14735_not n14736_not ; n14737
g14482 and b[6] n12668 ; n14738
g14483 and b[4] n13047 ; n14739
g14484 and b[5] n12663 ; n14740
g14485 and n14739_not n14740_not ; n14741
g14486 and n14738_not n14741 ; n14742
g14487 and n12671_not n14742 ; n14743
g14488 and n459_not n14742 ; n14744
g14489 and n14743_not n14744_not ; n14745
g14490 and a[62] n14745_not ; n14746
g14491 and a[62]_not n14745 ; n14747
g14492 and n14746_not n14747_not ; n14748
g14493 and n14737 n14748_not ; n14749
g14494 and n14737_not n14748 ; n14750
g14495 and n14749_not n14750_not ; n14751
g14496 and n14731_not n14751 ; n14752
g14497 and n14731 n14751_not ; n14753
g14498 and n14752_not n14753_not ; n14754
g14499 and b[9] n11531 ; n14755
g14500 and b[7] n11896 ; n14756
g14501 and b[8] n11526 ; n14757
g14502 and n14756_not n14757_not ; n14758
g14503 and n14755_not n14758 ; n14759
g14504 and n651 n11534 ; n14760
g14505 and n14759 n14760_not ; n14761
g14506 and a[59] n14761_not ; n14762
g14507 and a[59] n14762_not ; n14763
g14508 and n14761_not n14762_not ; n14764
g14509 and n14763_not n14764_not ; n14765
g14510 and n14754 n14765_not ; n14766
g14511 and n14754 n14766_not ; n14767
g14512 and n14765_not n14766_not ; n14768
g14513 and n14767_not n14768_not ; n14769
g14514 and n14275_not n14769 ; n14770
g14515 and n14275 n14769_not ; n14771
g14516 and n14770_not n14771_not ; n14772
g14517 and b[12] n10426 ; n14773
g14518 and b[10] n10796 ; n14774
g14519 and b[11] n10421 ; n14775
g14520 and n14774_not n14775_not ; n14776
g14521 and n14773_not n14776 ; n14777
g14522 and n842 n10429 ; n14778
g14523 and n14777 n14778_not ; n14779
g14524 and a[56] n14779_not ; n14780
g14525 and a[56] n14780_not ; n14781
g14526 and n14779_not n14780_not ; n14782
g14527 and n14781_not n14782_not ; n14783
g14528 and n14772 n14783 ; n14784
g14529 and n14772_not n14783_not ; n14785
g14530 and n14784_not n14785_not ; n14786
g14531 and n14730_not n14786 ; n14787
g14532 and n14730 n14786_not ; n14788
g14533 and n14787_not n14788_not ; n14789
g14534 and n14729_not n14789 ; n14790
g14535 and n14789 n14790_not ; n14791
g14536 and n14729_not n14790_not ; n14792
g14537 and n14791_not n14792_not ; n14793
g14538 and n14223_not n14298_not ; n14794
g14539 and n14295_not n14794_not ; n14795
g14540 and n14793 n14795 ; n14796
g14541 and n14793_not n14795_not ; n14797
g14542 and n14796_not n14797_not ; n14798
g14543 and b[18] n8362 ; n14799
g14544 and b[16] n8715 ; n14800
g14545 and b[17] n8357 ; n14801
g14546 and n14800_not n14801_not ; n14802
g14547 and n14799_not n14802 ; n14803
g14548 and n1566 n8365 ; n14804
g14549 and n14803 n14804_not ; n14805
g14550 and a[50] n14805_not ; n14806
g14551 and a[50] n14806_not ; n14807
g14552 and n14805_not n14806_not ; n14808
g14553 and n14807_not n14808_not ; n14809
g14554 and n14798 n14809_not ; n14810
g14555 and n14798 n14810_not ; n14811
g14556 and n14809_not n14810_not ; n14812
g14557 and n14811_not n14812_not ; n14813
g14558 and n14313_not n14317_not ; n14814
g14559 and n14813 n14814 ; n14815
g14560 and n14813_not n14814_not ; n14816
g14561 and n14815_not n14816_not ; n14817
g14562 and b[21] n7446 ; n14818
g14563 and b[19] n7787 ; n14819
g14564 and b[20] n7441 ; n14820
g14565 and n14819_not n14820_not ; n14821
g14566 and n14818_not n14821 ; n14822
g14567 and n1984 n7449 ; n14823
g14568 and n14822 n14823_not ; n14824
g14569 and a[47] n14824_not ; n14825
g14570 and a[47] n14825_not ; n14826
g14571 and n14824_not n14825_not ; n14827
g14572 and n14826_not n14827_not ; n14828
g14573 and n14817_not n14828 ; n14829
g14574 and n14817 n14828_not ; n14830
g14575 and n14829_not n14830_not ; n14831
g14576 and n14221_not n14333_not ; n14832
g14577 and n14330_not n14832_not ; n14833
g14578 and n14831 n14833_not ; n14834
g14579 and n14831_not n14833 ; n14835
g14580 and n14834_not n14835_not ; n14836
g14581 and n14718_not n14836 ; n14837
g14582 and n14836 n14837_not ; n14838
g14583 and n14718_not n14837_not ; n14839
g14584 and n14838_not n14839_not ; n14840
g14585 and n14348_not n14352_not ; n14841
g14586 and n14840 n14841 ; n14842
g14587 and n14840_not n14841_not ; n14843
g14588 and n14842_not n14843_not ; n14844
g14589 and b[27] n5777 ; n14845
g14590 and b[25] n6059 ; n14846
g14591 and b[26] n5772 ; n14847
g14592 and n14846_not n14847_not ; n14848
g14593 and n14845_not n14848 ; n14849
g14594 and n2990 n5780 ; n14850
g14595 and n14849 n14850_not ; n14851
g14596 and a[41] n14851_not ; n14852
g14597 and a[41] n14852_not ; n14853
g14598 and n14851_not n14852_not ; n14854
g14599 and n14853_not n14854_not ; n14855
g14600 and n14844 n14855_not ; n14856
g14601 and n14844 n14856_not ; n14857
g14602 and n14855_not n14856_not ; n14858
g14603 and n14857_not n14858_not ; n14859
g14604 and n14365_not n14371_not ; n14860
g14605 and n14859 n14860 ; n14861
g14606 and n14859_not n14860_not ; n14862
g14607 and n14861_not n14862_not ; n14863
g14608 and b[30] n5035 ; n14864
g14609 and b[28] n5277 ; n14865
g14610 and b[29] n5030 ; n14866
g14611 and n14865_not n14866_not ; n14867
g14612 and n14864_not n14867 ; n14868
g14613 and n3577 n5038 ; n14869
g14614 and n14868 n14869_not ; n14870
g14615 and a[38] n14870_not ; n14871
g14616 and a[38] n14871_not ; n14872
g14617 and n14870_not n14871_not ; n14873
g14618 and n14872_not n14873_not ; n14874
g14619 and n14863_not n14874 ; n14875
g14620 and n14863 n14874_not ; n14876
g14621 and n14875_not n14876_not ; n14877
g14622 and n14384_not n14390_not ; n14878
g14623 and n14877 n14878_not ; n14879
g14624 and n14877_not n14878 ; n14880
g14625 and n14879_not n14880_not ; n14881
g14626 and n14707_not n14881 ; n14882
g14627 and n14881 n14882_not ; n14883
g14628 and n14707_not n14882_not ; n14884
g14629 and n14883_not n14884_not ; n14885
g14630 and b[36] n3638 ; n14886
g14631 and b[34] n3843 ; n14887
g14632 and b[35] n3633 ; n14888
g14633 and n14887_not n14888_not ; n14889
g14634 and n14886_not n14889 ; n14890
g14635 and n3641_not n14890 ; n14891
g14636 and n4922_not n14890 ; n14892
g14637 and n14891_not n14892_not ; n14893
g14638 and a[32] n14893_not ; n14894
g14639 and a[32]_not n14893 ; n14895
g14640 and n14894_not n14895_not ; n14896
g14641 and n14408_not n14896_not ; n14897
g14642 and n14408_not n14897_not ; n14898
g14643 and n14896_not n14897_not ; n14899
g14644 and n14898_not n14899_not ; n14900
g14645 and n14885_not n14900_not ; n14901
g14646 and n14885_not n14901_not ; n14902
g14647 and n14900_not n14901_not ; n14903
g14648 and n14902_not n14903_not ; n14904
g14649 and n14696 n14904_not ; n14905
g14650 and n14696 n14905_not ; n14906
g14651 and n14904_not n14905_not ; n14907
g14652 and n14906_not n14907_not ; n14908
g14653 and n14681 n14908_not ; n14909
g14654 and n14681_not n14908 ; n14910
g14655 and n14666_not n14910_not ; n14911
g14656 and n14909_not n14911 ; n14912
g14657 and n14666_not n14912_not ; n14913
g14658 and n14910_not n14912_not ; n14914
g14659 and n14909_not n14914 ; n14915
g14660 and n14913_not n14915_not ; n14916
g14661 and n14652 n14916_not ; n14917
g14662 and n14652_not n14916 ; n14918
g14663 and n14637 n14918_not ; n14919
g14664 and n14917_not n14919 ; n14920
g14665 and n14637 n14920_not ; n14921
g14666 and n14918_not n14920_not ; n14922
g14667 and n14917_not n14922 ; n14923
g14668 and n14921_not n14923_not ; n14924
g14669 and n14508_not n14510_not ; n14925
g14670 and b[54] n951 ; n14926
g14671 and b[52] n1056 ; n14927
g14672 and b[53] n946 ; n14928
g14673 and n14927_not n14928_not ; n14929
g14674 and n14926_not n14929 ; n14930
g14675 and n954_not n14930 ; n14931
g14676 and n9998_not n14930 ; n14932
g14677 and n14931_not n14932_not ; n14933
g14678 and a[14] n14933_not ; n14934
g14679 and a[14]_not n14933 ; n14935
g14680 and n14934_not n14935_not ; n14936
g14681 and n14925_not n14936_not ; n14937
g14682 and n14925_not n14937_not ; n14938
g14683 and n14936_not n14937_not ; n14939
g14684 and n14938_not n14939_not ; n14940
g14685 and n14924_not n14940_not ; n14941
g14686 and n14924_not n14941_not ; n14942
g14687 and n14940_not n14941_not ; n14943
g14688 and n14942_not n14943_not ; n14944
g14689 and n14622 n14944_not ; n14945
g14690 and n14622 n14945_not ; n14946
g14691 and n14944_not n14945_not ; n14947
g14692 and n14946_not n14947_not ; n14948
g14693 and b[60] n511 ; n14949
g14694 and b[58] n541 ; n14950
g14695 and b[59] n506 ; n14951
g14696 and n14950_not n14951_not ; n14952
g14697 and n14949_not n14952 ; n14953
g14698 and n514 n12211 ; n14954
g14699 and n14953 n14954_not ; n14955
g14700 and a[8] n14955_not ; n14956
g14701 and a[8] n14956_not ; n14957
g14702 and n14955_not n14956_not ; n14958
g14703 and n14957_not n14958_not ; n14959
g14704 and n14533_not n14546_not ; n14960
g14705 and n14959_not n14960_not ; n14961
g14706 and n14959_not n14961_not ; n14962
g14707 and n14960_not n14961_not ; n14963
g14708 and n14962_not n14963_not ; n14964
g14709 and n14948_not n14964_not ; n14965
g14710 and n14948_not n14965_not ; n14966
g14711 and n14964_not n14965_not ; n14967
g14712 and n14966_not n14967_not ; n14968
g14713 and n14607_not n14968_not ; n14969
g14714 and n14607_not n14969_not ; n14970
g14715 and n14968_not n14969_not ; n14971
g14716 and n14970_not n14971_not ; n14972
g14717 and n14577_not n14580_not ; n14973
g14718 and n14972 n14973 ; n14974
g14719 and n14972_not n14973_not ; n14975
g14720 and n14974_not n14975_not ; n14976
g14721 and n14586_not n14589_not ; n14977
g14722 and n14976 n14977_not ; n14978
g14723 and n14976_not n14977 ; n14979
g14724 and n14978_not n14979_not ; f[66]
g14725 and n14975_not n14978_not ; n14981
g14726 and n14604_not n14969_not ; n14982
g14727 and b[55] n951 ; n14983
g14728 and b[53] n1056 ; n14984
g14729 and b[54] n946 ; n14985
g14730 and n14984_not n14985_not ; n14986
g14731 and n14983_not n14986 ; n14987
g14732 and n954 n10684 ; n14988
g14733 and n14987 n14988_not ; n14989
g14734 and a[14] n14989_not ; n14990
g14735 and a[14] n14990_not ; n14991
g14736 and n14989_not n14990_not ; n14992
g14737 and n14991_not n14992_not ; n14993
g14738 and n14636_not n14920_not ; n14994
g14739 and n14993 n14994 ; n14995
g14740 and n14993_not n14994_not ; n14996
g14741 and n14995_not n14996_not ; n14997
g14742 and b[49] n1627 ; n14998
g14743 and b[47] n1763 ; n14999
g14744 and b[48] n1622 ; n15000
g14745 and n14999_not n15000_not ; n15001
g14746 and n14998_not n15001 ; n15002
g14747 and n1630 n8625 ; n15003
g14748 and n15002 n15003_not ; n15004
g14749 and a[20] n15004_not ; n15005
g14750 and a[20] n15005_not ; n15006
g14751 and n15004_not n15005_not ; n15007
g14752 and n15006_not n15007_not ; n15008
g14753 and n14465_not n14663_not ; n15009
g14754 and n14912_not n15009_not ; n15010
g14755 and n15008 n15010 ; n15011
g14756 and n15008_not n15010_not ; n15012
g14757 and n15011_not n15012_not ; n15013
g14758 and b[43] n2539 ; n15014
g14759 and b[41] n2685 ; n15015
g14760 and b[42] n2534 ; n15016
g14761 and n15015_not n15016_not ; n15017
g14762 and n15014_not n15017 ; n15018
g14763 and n2542 n6515 ; n15019
g14764 and n15018 n15019_not ; n15020
g14765 and a[26] n15020_not ; n15021
g14766 and a[26] n15021_not ; n15022
g14767 and n15020_not n15021_not ; n15023
g14768 and n15022_not n15023_not ; n15024
g14769 and n14694_not n14905_not ; n15025
g14770 and n15024 n15025 ; n15026
g14771 and n15024_not n15025_not ; n15027
g14772 and n15026_not n15027_not ; n15028
g14773 and n14879_not n14882_not ; n15029
g14774 and b[37] n3638 ; n15030
g14775 and b[35] n3843 ; n15031
g14776 and b[36] n3633 ; n15032
g14777 and n15031_not n15032_not ; n15033
g14778 and n15030_not n15033 ; n15034
g14779 and n3641_not n15034 ; n15035
g14780 and n5181_not n15034 ; n15036
g14781 and n15035_not n15036_not ; n15037
g14782 and a[32] n15037_not ; n15038
g14783 and a[32]_not n15037 ; n15039
g14784 and n15038_not n15039_not ; n15040
g14785 and n15029_not n15040_not ; n15041
g14786 and n15029 n15040 ; n15042
g14787 and n15041_not n15042_not ; n15043
g14788 and b[34] n4287 ; n15044
g14789 and b[32] n4532 ; n15045
g14790 and b[33] n4282 ; n15046
g14791 and n15045_not n15046_not ; n15047
g14792 and n15044_not n15047 ; n15048
g14793 and n4290 n4466 ; n15049
g14794 and n15048 n15049_not ; n15050
g14795 and a[35] n15050_not ; n15051
g14796 and a[35] n15051_not ; n15052
g14797 and n15050_not n15051_not ; n15053
g14798 and n15052_not n15053_not ; n15054
g14799 and n14862_not n14876_not ; n15055
g14800 and b[16] n9339 ; n15056
g14801 and b[14] n9732 ; n15057
g14802 and b[15] n9334 ; n15058
g14803 and n15057_not n15058_not ; n15059
g14804 and n15056_not n15059 ; n15060
g14805 and n1237 n9342 ; n15061
g14806 and n15060 n15061_not ; n15062
g14807 and a[53] n15062_not ; n15063
g14808 and a[53] n15063_not ; n15064
g14809 and n15062_not n15063_not ; n15065
g14810 and n15064_not n15065_not ; n15066
g14811 and b[7] n12668 ; n15067
g14812 and b[5] n13047 ; n15068
g14813 and b[6] n12663 ; n15069
g14814 and n15068_not n15069_not ; n15070
g14815 and n15067_not n15070 ; n15071
g14816 and n484 n12671 ; n15072
g14817 and n15071 n15072_not ; n15073
g14818 and a[62] n15073_not ; n15074
g14819 and a[62] n15074_not ; n15075
g14820 and n15073_not n15074_not ; n15076
g14821 and n15075_not n15076_not ; n15077
g14822 and b[3] n13903 ; n15078
g14823 and b[4] n13488_not ; n15079
g14824 and n15078_not n15079_not ; n15080
g14825 and a[2] n15080_not ; n15081
g14826 and a[2] n15081_not ; n15082
g14827 and n15080_not n15081_not ; n15083
g14828 and n15082_not n15083_not ; n15084
g14829 and n15077_not n15084_not ; n15085
g14830 and n15077_not n15085_not ; n15086
g14831 and n15084_not n15085_not ; n15087
g14832 and n15086_not n15087_not ; n15088
g14833 and n14735_not n14749_not ; n15089
g14834 and n15088 n15089 ; n15090
g14835 and n15088_not n15089_not ; n15091
g14836 and n15090_not n15091_not ; n15092
g14837 and b[10] n11531 ; n15093
g14838 and b[8] n11896 ; n15094
g14839 and b[9] n11526 ; n15095
g14840 and n15094_not n15095_not ; n15096
g14841 and n15093_not n15096 ; n15097
g14842 and n738 n11534 ; n15098
g14843 and n15097 n15098_not ; n15099
g14844 and a[59] n15099_not ; n15100
g14845 and a[59] n15100_not ; n15101
g14846 and n15099_not n15100_not ; n15102
g14847 and n15101_not n15102_not ; n15103
g14848 and n15092 n15103_not ; n15104
g14849 and n15092 n15104_not ; n15105
g14850 and n15103_not n15104_not ; n15106
g14851 and n15105_not n15106_not ; n15107
g14852 and n14752_not n14766_not ; n15108
g14853 and n15107 n15108 ; n15109
g14854 and n15107_not n15108_not ; n15110
g14855 and n15109_not n15110_not ; n15111
g14856 and b[13] n10426 ; n15112
g14857 and b[11] n10796 ; n15113
g14858 and b[12] n10421 ; n15114
g14859 and n15113_not n15114_not ; n15115
g14860 and n15112_not n15115 ; n15116
g14861 and n1008 n10429 ; n15117
g14862 and n15116 n15117_not ; n15118
g14863 and a[56] n15118_not ; n15119
g14864 and a[56] n15119_not ; n15120
g14865 and n15118_not n15119_not ; n15121
g14866 and n15120_not n15121_not ; n15122
g14867 and n15111_not n15122 ; n15123
g14868 and n15111 n15122_not ; n15124
g14869 and n15123_not n15124_not ; n15125
g14870 and n14275_not n14769_not ; n15126
g14871 and n14785_not n15126_not ; n15127
g14872 and n15125 n15127_not ; n15128
g14873 and n15125_not n15127 ; n15129
g14874 and n15128_not n15129_not ; n15130
g14875 and n15066_not n15130 ; n15131
g14876 and n15130 n15131_not ; n15132
g14877 and n15066_not n15131_not ; n15133
g14878 and n15132_not n15133_not ; n15134
g14879 and n14787_not n14790_not ; n15135
g14880 and n15134 n15135 ; n15136
g14881 and n15134_not n15135_not ; n15137
g14882 and n15136_not n15137_not ; n15138
g14883 and b[19] n8362 ; n15139
g14884 and b[17] n8715 ; n15140
g14885 and b[18] n8357 ; n15141
g14886 and n15140_not n15141_not ; n15142
g14887 and n15139_not n15142 ; n15143
g14888 and n1708 n8365 ; n15144
g14889 and n15143 n15144_not ; n15145
g14890 and a[50] n15145_not ; n15146
g14891 and a[50] n15146_not ; n15147
g14892 and n15145_not n15146_not ; n15148
g14893 and n15147_not n15148_not ; n15149
g14894 and n15138 n15149_not ; n15150
g14895 and n15138 n15150_not ; n15151
g14896 and n15149_not n15150_not ; n15152
g14897 and n15151_not n15152_not ; n15153
g14898 and n14797_not n14810_not ; n15154
g14899 and n15153 n15154 ; n15155
g14900 and n15153_not n15154_not ; n15156
g14901 and n15155_not n15156_not ; n15157
g14902 and b[22] n7446 ; n15158
g14903 and b[20] n7787 ; n15159
g14904 and b[21] n7441 ; n15160
g14905 and n15159_not n15160_not ; n15161
g14906 and n15158_not n15161 ; n15162
g14907 and n2145 n7449 ; n15163
g14908 and n15162 n15163_not ; n15164
g14909 and a[47] n15164_not ; n15165
g14910 and a[47] n15165_not ; n15166
g14911 and n15164_not n15165_not ; n15167
g14912 and n15166_not n15167_not ; n15168
g14913 and n15157 n15168_not ; n15169
g14914 and n15157 n15169_not ; n15170
g14915 and n15168_not n15169_not ; n15171
g14916 and n15170_not n15171_not ; n15172
g14917 and n14816_not n14830_not ; n15173
g14918 and n15172_not n15173_not ; n15174
g14919 and n15172_not n15174_not ; n15175
g14920 and n15173_not n15174_not ; n15176
g14921 and n15175_not n15176_not ; n15177
g14922 and b[25] n6595 ; n15178
g14923 and b[23] n6902 ; n15179
g14924 and b[24] n6590 ; n15180
g14925 and n15179_not n15180_not ; n15181
g14926 and n15178_not n15181 ; n15182
g14927 and n2485 n6598 ; n15183
g14928 and n15182 n15183_not ; n15184
g14929 and a[44] n15184_not ; n15185
g14930 and a[44] n15185_not ; n15186
g14931 and n15184_not n15185_not ; n15187
g14932 and n15186_not n15187_not ; n15188
g14933 and n15177_not n15188_not ; n15189
g14934 and n15177_not n15189_not ; n15190
g14935 and n15188_not n15189_not ; n15191
g14936 and n15190_not n15191_not ; n15192
g14937 and n14834_not n14837_not ; n15193
g14938 and n15192 n15193 ; n15194
g14939 and n15192_not n15193_not ; n15195
g14940 and n15194_not n15195_not ; n15196
g14941 and b[28] n5777 ; n15197
g14942 and b[26] n6059 ; n15198
g14943 and b[27] n5772 ; n15199
g14944 and n15198_not n15199_not ; n15200
g14945 and n15197_not n15200 ; n15201
g14946 and n3189 n5780 ; n15202
g14947 and n15201 n15202_not ; n15203
g14948 and a[41] n15203_not ; n15204
g14949 and a[41] n15204_not ; n15205
g14950 and n15203_not n15204_not ; n15206
g14951 and n15205_not n15206_not ; n15207
g14952 and n15196 n15207_not ; n15208
g14953 and n15196 n15208_not ; n15209
g14954 and n15207_not n15208_not ; n15210
g14955 and n15209_not n15210_not ; n15211
g14956 and n14843_not n14856_not ; n15212
g14957 and n15211 n15212 ; n15213
g14958 and n15211_not n15212_not ; n15214
g14959 and n15213_not n15214_not ; n15215
g14960 and b[31] n5035 ; n15216
g14961 and b[29] n5277 ; n15217
g14962 and b[30] n5030 ; n15218
g14963 and n15217_not n15218_not ; n15219
g14964 and n15216_not n15219 ; n15220
g14965 and n3796 n5038 ; n15221
g14966 and n15220 n15221_not ; n15222
g14967 and a[38] n15222_not ; n15223
g14968 and a[38] n15223_not ; n15224
g14969 and n15222_not n15223_not ; n15225
g14970 and n15224_not n15225_not ; n15226
g14971 and n15215_not n15226 ; n15227
g14972 and n15215 n15226_not ; n15228
g14973 and n15227_not n15228_not ; n15229
g14974 and n15055_not n15229 ; n15230
g14975 and n15055_not n15230_not ; n15231
g14976 and n15229 n15230_not ; n15232
g14977 and n15231_not n15232_not ; n15233
g14978 and n15054_not n15233_not ; n15234
g14979 and n15054_not n15234_not ; n15235
g14980 and n15233_not n15234_not ; n15236
g14981 and n15235_not n15236_not ; n15237
g14982 and n15043_not n15237 ; n15238
g14983 and n15043 n15237_not ; n15239
g14984 and n15238_not n15239_not ; n15240
g14985 and n14897_not n14901_not ; n15241
g14986 and b[40] n3050 ; n15242
g14987 and b[38] n3243 ; n15243
g14988 and b[39] n3045 ; n15244
g14989 and n15243_not n15244_not ; n15245
g14990 and n15242_not n15245 ; n15246
g14991 and n3053_not n15246 ; n15247
g14992 and n5955_not n15246 ; n15248
g14993 and n15247_not n15248_not ; n15249
g14994 and a[29] n15249_not ; n15250
g14995 and a[29]_not n15249 ; n15251
g14996 and n15250_not n15251_not ; n15252
g14997 and n15241_not n15252_not ; n15253
g14998 and n15241_not n15253_not ; n15254
g14999 and n15252_not n15253_not ; n15255
g15000 and n15254_not n15255_not ; n15256
g15001 and n15240 n15256_not ; n15257
g15002 and n15240 n15257_not ; n15258
g15003 and n15256_not n15257_not ; n15259
g15004 and n15258_not n15259_not ; n15260
g15005 and n15028 n15260_not ; n15261
g15006 and n15028 n15261_not ; n15262
g15007 and n15260_not n15261_not ; n15263
g15008 and n15262_not n15263_not ; n15264
g15009 and b[46] n2048 ; n15265
g15010 and b[44] n2198 ; n15266
g15011 and b[45] n2043 ; n15267
g15012 and n15266_not n15267_not ; n15268
g15013 and n15265_not n15268 ; n15269
g15014 and n2051 n7677 ; n15270
g15015 and n15269 n15270_not ; n15271
g15016 and a[23] n15271_not ; n15272
g15017 and a[23] n15272_not ; n15273
g15018 and n15271_not n15272_not ; n15274
g15019 and n15273_not n15274_not ; n15275
g15020 and n14680_not n14909_not ; n15276
g15021 and n15275_not n15276_not ; n15277
g15022 and n15275_not n15277_not ; n15278
g15023 and n15276_not n15277_not ; n15279
g15024 and n15278_not n15279_not ; n15280
g15025 and n15264_not n15280 ; n15281
g15026 and n15264 n15280_not ; n15282
g15027 and n15281_not n15282_not ; n15283
g15028 and n15013 n15283_not ; n15284
g15029 and n15013 n15284_not ; n15285
g15030 and n15283_not n15284_not ; n15286
g15031 and n15285_not n15286_not ; n15287
g15032 and b[52] n1302 ; n15288
g15033 and b[50] n1391 ; n15289
g15034 and b[51] n1297 ; n15290
g15035 and n15289_not n15290_not ; n15291
g15036 and n15288_not n15291 ; n15292
g15037 and n1305 n9628 ; n15293
g15038 and n15292 n15293_not ; n15294
g15039 and a[17] n15294_not ; n15295
g15040 and a[17] n15295_not ; n15296
g15041 and n15294_not n15295_not ; n15297
g15042 and n15296_not n15297_not ; n15298
g15043 and n14651_not n14917_not ; n15299
g15044 and n15298_not n15299_not ; n15300
g15045 and n15298_not n15300_not ; n15301
g15046 and n15299_not n15300_not ; n15302
g15047 and n15301_not n15302_not ; n15303
g15048 and n15287_not n15303 ; n15304
g15049 and n15287 n15303_not ; n15305
g15050 and n15304_not n15305_not ; n15306
g15051 and n14997 n15306_not ; n15307
g15052 and n14997 n15307_not ; n15308
g15053 and n15306_not n15307_not ; n15309
g15054 and n15308_not n15309_not ; n15310
g15055 and n14937_not n14941_not ; n15311
g15056 and b[58] n700 ; n15312
g15057 and b[56] n767 ; n15313
g15058 and b[57] n695 ; n15314
g15059 and n15313_not n15314_not ; n15315
g15060 and n15312_not n15315 ; n15316
g15061 and n703_not n15316 ; n15317
g15062 and n11436_not n15316 ; n15318
g15063 and n15317_not n15318_not ; n15319
g15064 and a[11] n15319_not ; n15320
g15065 and a[11]_not n15319 ; n15321
g15066 and n15320_not n15321_not ; n15322
g15067 and n15311_not n15322_not ; n15323
g15068 and n15311_not n15323_not ; n15324
g15069 and n15322_not n15323_not ; n15325
g15070 and n15324_not n15325_not ; n15326
g15071 and n15310_not n15326_not ; n15327
g15072 and n15310_not n15327_not ; n15328
g15073 and n15326_not n15327_not ; n15329
g15074 and n15328_not n15329_not ; n15330
g15075 and n14621_not n14945_not ; n15331
g15076 and b[61] n511 ; n15332
g15077 and b[59] n541 ; n15333
g15078 and b[60] n506 ; n15334
g15079 and n15333_not n15334_not ; n15335
g15080 and n15332_not n15335 ; n15336
g15081 and n514_not n15336 ; n15337
g15082 and n12969_not n15336 ; n15338
g15083 and n15337_not n15338_not ; n15339
g15084 and a[8] n15339_not ; n15340
g15085 and a[8]_not n15339 ; n15341
g15086 and n15340_not n15341_not ; n15342
g15087 and n15331_not n15342_not ; n15343
g15088 and n15331_not n15343_not ; n15344
g15089 and n15342_not n15343_not ; n15345
g15090 and n15344_not n15345_not ; n15346
g15091 and n15330_not n15346_not ; n15347
g15092 and n15330_not n15347_not ; n15348
g15093 and n15346_not n15347_not ; n15349
g15094 and n15348_not n15349_not ; n15350
g15095 and n14961_not n14965_not ; n15351
g15096 and b[62] n403 ; n15352
g15097 and b[63] n357 ; n15353
g15098 and n15352_not n15353_not ; n15354
g15099 and n365_not n15354 ; n15355
g15100 and n13800 n15354 ; n15356
g15101 and n15355_not n15356_not ; n15357
g15102 and a[5] n15357_not ; n15358
g15103 and a[5]_not n15357 ; n15359
g15104 and n15358_not n15359_not ; n15360
g15105 and n15351_not n15360_not ; n15361
g15106 and n15351_not n15361_not ; n15362
g15107 and n15360_not n15361_not ; n15363
g15108 and n15362_not n15363_not ; n15364
g15109 and n15350_not n15364_not ; n15365
g15110 and n15350 n15363_not ; n15366
g15111 and n15362_not n15366 ; n15367
g15112 and n15365_not n15367_not ; n15368
g15113 and n14982_not n15368 ; n15369
g15114 and n14982_not n15369_not ; n15370
g15115 and n15368 n15369_not ; n15371
g15116 and n15370_not n15371_not ; n15372
g15117 and n14981_not n15372_not ; n15373
g15118 and n14981 n15371_not ; n15374
g15119 and n15370_not n15374 ; n15375
g15120 and n15373_not n15375_not ; f[67]
g15121 and n15369_not n15373_not ; n15377
g15122 and n15361_not n15365_not ; n15378
g15123 and n15343_not n15347_not ; n15379
g15124 and b[63] n403 ; n15380
g15125 and n365 n13797 ; n15381
g15126 and n15380_not n15381_not ; n15382
g15127 and a[5] n15382_not ; n15383
g15128 and a[5] n15383_not ; n15384
g15129 and n15382_not n15383_not ; n15385
g15130 and n15384_not n15385_not ; n15386
g15131 and n15379_not n15386_not ; n15387
g15132 and n15379_not n15387_not ; n15388
g15133 and n15386_not n15387_not ; n15389
g15134 and n15388_not n15389_not ; n15390
g15135 and b[59] n700 ; n15391
g15136 and b[57] n767 ; n15392
g15137 and b[58] n695 ; n15393
g15138 and n15392_not n15393_not ; n15394
g15139 and n15391_not n15394 ; n15395
g15140 and n703 n12179 ; n15396
g15141 and n15395 n15396_not ; n15397
g15142 and a[11] n15397_not ; n15398
g15143 and a[11] n15398_not ; n15399
g15144 and n15397_not n15398_not ; n15400
g15145 and n15399_not n15400_not ; n15401
g15146 and n14996_not n15307_not ; n15402
g15147 and n15401 n15402 ; n15403
g15148 and n15401_not n15402_not ; n15404
g15149 and n15403_not n15404_not ; n15405
g15150 and b[56] n951 ; n15406
g15151 and b[54] n1056 ; n15407
g15152 and b[55] n946 ; n15408
g15153 and n15407_not n15408_not ; n15409
g15154 and n15406_not n15409 ; n15410
g15155 and n954 n10708 ; n15411
g15156 and n15410 n15411_not ; n15412
g15157 and a[14] n15412_not ; n15413
g15158 and a[14] n15413_not ; n15414
g15159 and n15412_not n15413_not ; n15415
g15160 and n15414_not n15415_not ; n15416
g15161 and n15287_not n15303_not ; n15417
g15162 and n15300_not n15417_not ; n15418
g15163 and n15416_not n15418_not ; n15419
g15164 and n15416_not n15419_not ; n15420
g15165 and n15418_not n15419_not ; n15421
g15166 and n15420_not n15421_not ; n15422
g15167 and n15012_not n15284_not ; n15423
g15168 and b[53] n1302 ; n15424
g15169 and b[51] n1391 ; n15425
g15170 and b[52] n1297 ; n15426
g15171 and n15425_not n15426_not ; n15427
g15172 and n15424_not n15427 ; n15428
g15173 and n1305_not n15428 ; n15429
g15174 and n9972_not n15428 ; n15430
g15175 and n15429_not n15430_not ; n15431
g15176 and a[17] n15431_not ; n15432
g15177 and a[17]_not n15431 ; n15433
g15178 and n15432_not n15433_not ; n15434
g15179 and n15423_not n15434_not ; n15435
g15180 and n15423 n15434 ; n15436
g15181 and n15435_not n15436_not ; n15437
g15182 and b[50] n1627 ; n15438
g15183 and b[48] n1763 ; n15439
g15184 and b[49] n1622 ; n15440
g15185 and n15439_not n15440_not ; n15441
g15186 and n15438_not n15441 ; n15442
g15187 and n1630 n8949 ; n15443
g15188 and n15442 n15443_not ; n15444
g15189 and a[20] n15444_not ; n15445
g15190 and a[20] n15445_not ; n15446
g15191 and n15444_not n15445_not ; n15447
g15192 and n15446_not n15447_not ; n15448
g15193 and n15264_not n15280_not ; n15449
g15194 and n15277_not n15449_not ; n15450
g15195 and n15448_not n15450_not ; n15451
g15196 and n15448_not n15451_not ; n15452
g15197 and n15450_not n15451_not ; n15453
g15198 and n15452_not n15453_not ; n15454
g15199 and b[47] n2048 ; n15455
g15200 and b[45] n2198 ; n15456
g15201 and b[46] n2043 ; n15457
g15202 and n15456_not n15457_not ; n15458
g15203 and n15455_not n15458 ; n15459
g15204 and n2051 n7703 ; n15460
g15205 and n15459 n15460_not ; n15461
g15206 and a[23] n15461_not ; n15462
g15207 and a[23] n15462_not ; n15463
g15208 and n15461_not n15462_not ; n15464
g15209 and n15463_not n15464_not ; n15465
g15210 and n15027_not n15261_not ; n15466
g15211 and n15465 n15466 ; n15467
g15212 and n15465_not n15466_not ; n15468
g15213 and n15467_not n15468_not ; n15469
g15214 and b[41] n3050 ; n15470
g15215 and b[39] n3243 ; n15471
g15216 and b[40] n3045 ; n15472
g15217 and n15471_not n15472_not ; n15473
g15218 and n15470_not n15473 ; n15474
g15219 and n3053 n6219 ; n15475
g15220 and n15474 n15475_not ; n15476
g15221 and a[29] n15476_not ; n15477
g15222 and a[29] n15477_not ; n15478
g15223 and n15476_not n15477_not ; n15479
g15224 and n15478_not n15479_not ; n15480
g15225 and n15041_not n15239_not ; n15481
g15226 and n15480 n15481 ; n15482
g15227 and n15480_not n15481_not ; n15483
g15228 and n15482_not n15483_not ; n15484
g15229 and b[35] n4287 ; n15485
g15230 and b[33] n4532 ; n15486
g15231 and b[34] n4282 ; n15487
g15232 and n15486_not n15487_not ; n15488
g15233 and n15485_not n15488 ; n15489
g15234 and n4290 n4696 ; n15490
g15235 and n15489 n15490_not ; n15491
g15236 and a[35] n15491_not ; n15492
g15237 and a[35] n15492_not ; n15493
g15238 and n15491_not n15492_not ; n15494
g15239 and n15493_not n15494_not ; n15495
g15240 and b[23] n7446 ; n15496
g15241 and b[21] n7787 ; n15497
g15242 and b[22] n7441 ; n15498
g15243 and n15497_not n15498_not ; n15499
g15244 and n15496_not n15499 ; n15500
g15245 and n2300 n7449 ; n15501
g15246 and n15500 n15501_not ; n15502
g15247 and a[47] n15502_not ; n15503
g15248 and a[47] n15503_not ; n15504
g15249 and n15502_not n15503_not ; n15505
g15250 and n15504_not n15505_not ; n15506
g15251 and b[14] n10426 ; n15507
g15252 and b[12] n10796 ; n15508
g15253 and b[13] n10421 ; n15509
g15254 and n15508_not n15509_not ; n15510
g15255 and n15507_not n15510 ; n15511
g15256 and n1034 n10429 ; n15512
g15257 and n15511 n15512_not ; n15513
g15258 and a[56] n15513_not ; n15514
g15259 and a[56] n15514_not ; n15515
g15260 and n15513_not n15514_not ; n15516
g15261 and n15515_not n15516_not ; n15517
g15262 and b[8] n12668 ; n15518
g15263 and b[6] n13047 ; n15519
g15264 and b[7] n12663 ; n15520
g15265 and n15519_not n15520_not ; n15521
g15266 and n15518_not n15521 ; n15522
g15267 and n585 n12671 ; n15523
g15268 and n15522 n15523_not ; n15524
g15269 and a[62] n15524_not ; n15525
g15270 and a[62] n15525_not ; n15526
g15271 and n15524_not n15525_not ; n15527
g15272 and n15526_not n15527_not ; n15528
g15273 and b[4] n13903 ; n15529
g15274 and b[5] n13488_not ; n15530
g15275 and n15529_not n15530_not ; n15531
g15276 and a[2] n15531_not ; n15532
g15277 and a[2] n15532_not ; n15533
g15278 and n15531_not n15532_not ; n15534
g15279 and n15533_not n15534_not ; n15535
g15280 and n15528_not n15535_not ; n15536
g15281 and n15528_not n15536_not ; n15537
g15282 and n15535_not n15536_not ; n15538
g15283 and n15537_not n15538_not ; n15539
g15284 and n15081_not n15085_not ; n15540
g15285 and n15539 n15540 ; n15541
g15286 and n15539_not n15540_not ; n15542
g15287 and n15541_not n15542_not ; n15543
g15288 and b[11] n11531 ; n15544
g15289 and b[9] n11896 ; n15545
g15290 and b[10] n11526 ; n15546
g15291 and n15545_not n15546_not ; n15547
g15292 and n15544_not n15547 ; n15548
g15293 and n818 n11534 ; n15549
g15294 and n15548 n15549_not ; n15550
g15295 and a[59] n15550_not ; n15551
g15296 and a[59] n15551_not ; n15552
g15297 and n15550_not n15551_not ; n15553
g15298 and n15552_not n15553_not ; n15554
g15299 and n15543_not n15554 ; n15555
g15300 and n15543 n15554_not ; n15556
g15301 and n15555_not n15556_not ; n15557
g15302 and n15091_not n15104_not ; n15558
g15303 and n15557 n15558_not ; n15559
g15304 and n15557_not n15558 ; n15560
g15305 and n15559_not n15560_not ; n15561
g15306 and n15517_not n15561 ; n15562
g15307 and n15561 n15562_not ; n15563
g15308 and n15517_not n15562_not ; n15564
g15309 and n15563_not n15564_not ; n15565
g15310 and n15110_not n15124_not ; n15566
g15311 and n15565_not n15566_not ; n15567
g15312 and n15565_not n15567_not ; n15568
g15313 and n15566_not n15567_not ; n15569
g15314 and n15568_not n15569_not ; n15570
g15315 and b[17] n9339 ; n15571
g15316 and b[15] n9732 ; n15572
g15317 and b[16] n9334 ; n15573
g15318 and n15572_not n15573_not ; n15574
g15319 and n15571_not n15574 ; n15575
g15320 and n1356 n9342 ; n15576
g15321 and n15575 n15576_not ; n15577
g15322 and a[53] n15577_not ; n15578
g15323 and a[53] n15578_not ; n15579
g15324 and n15577_not n15578_not ; n15580
g15325 and n15579_not n15580_not ; n15581
g15326 and n15570_not n15581_not ; n15582
g15327 and n15570_not n15582_not ; n15583
g15328 and n15581_not n15582_not ; n15584
g15329 and n15583_not n15584_not ; n15585
g15330 and n15128_not n15131_not ; n15586
g15331 and n15585 n15586 ; n15587
g15332 and n15585_not n15586_not ; n15588
g15333 and n15587_not n15588_not ; n15589
g15334 and b[20] n8362 ; n15590
g15335 and b[18] n8715 ; n15591
g15336 and b[19] n8357 ; n15592
g15337 and n15591_not n15592_not ; n15593
g15338 and n15590_not n15593 ; n15594
g15339 and n1846 n8365 ; n15595
g15340 and n15594 n15595_not ; n15596
g15341 and a[50] n15596_not ; n15597
g15342 and a[50] n15597_not ; n15598
g15343 and n15596_not n15597_not ; n15599
g15344 and n15598_not n15599_not ; n15600
g15345 and n15589_not n15600 ; n15601
g15346 and n15589 n15600_not ; n15602
g15347 and n15601_not n15602_not ; n15603
g15348 and n15137_not n15150_not ; n15604
g15349 and n15603 n15604_not ; n15605
g15350 and n15603_not n15604 ; n15606
g15351 and n15605_not n15606_not ; n15607
g15352 and n15506_not n15607 ; n15608
g15353 and n15607 n15608_not ; n15609
g15354 and n15506_not n15608_not ; n15610
g15355 and n15609_not n15610_not ; n15611
g15356 and n15156_not n15169_not ; n15612
g15357 and n15611 n15612 ; n15613
g15358 and n15611_not n15612_not ; n15614
g15359 and n15613_not n15614_not ; n15615
g15360 and b[26] n6595 ; n15616
g15361 and b[24] n6902 ; n15617
g15362 and b[25] n6590 ; n15618
g15363 and n15617_not n15618_not ; n15619
g15364 and n15616_not n15619 ; n15620
g15365 and n2813 n6598 ; n15621
g15366 and n15620 n15621_not ; n15622
g15367 and a[44] n15622_not ; n15623
g15368 and a[44] n15623_not ; n15624
g15369 and n15622_not n15623_not ; n15625
g15370 and n15624_not n15625_not ; n15626
g15371 and n15615 n15626_not ; n15627
g15372 and n15615 n15627_not ; n15628
g15373 and n15626_not n15627_not ; n15629
g15374 and n15628_not n15629_not ; n15630
g15375 and n15174_not n15189_not ; n15631
g15376 and n15630 n15631 ; n15632
g15377 and n15630_not n15631_not ; n15633
g15378 and n15632_not n15633_not ; n15634
g15379 and b[29] n5777 ; n15635
g15380 and b[27] n6059 ; n15636
g15381 and b[28] n5772 ; n15637
g15382 and n15636_not n15637_not ; n15638
g15383 and n15635_not n15638 ; n15639
g15384 and n3383 n5780 ; n15640
g15385 and n15639 n15640_not ; n15641
g15386 and a[41] n15641_not ; n15642
g15387 and a[41] n15642_not ; n15643
g15388 and n15641_not n15642_not ; n15644
g15389 and n15643_not n15644_not ; n15645
g15390 and n15634 n15645_not ; n15646
g15391 and n15634 n15646_not ; n15647
g15392 and n15645_not n15646_not ; n15648
g15393 and n15647_not n15648_not ; n15649
g15394 and n15195_not n15208_not ; n15650
g15395 and n15649 n15650 ; n15651
g15396 and n15649_not n15650_not ; n15652
g15397 and n15651_not n15652_not ; n15653
g15398 and b[32] n5035 ; n15654
g15399 and b[30] n5277 ; n15655
g15400 and b[31] n5030 ; n15656
g15401 and n15655_not n15656_not ; n15657
g15402 and n15654_not n15657 ; n15658
g15403 and n4013 n5038 ; n15659
g15404 and n15658 n15659_not ; n15660
g15405 and a[38] n15660_not ; n15661
g15406 and a[38] n15661_not ; n15662
g15407 and n15660_not n15661_not ; n15663
g15408 and n15662_not n15663_not ; n15664
g15409 and n15653_not n15664 ; n15665
g15410 and n15653 n15664_not ; n15666
g15411 and n15665_not n15666_not ; n15667
g15412 and n15214_not n15228_not ; n15668
g15413 and n15667 n15668_not ; n15669
g15414 and n15667_not n15668 ; n15670
g15415 and n15669_not n15670_not ; n15671
g15416 and n15495_not n15671 ; n15672
g15417 and n15671 n15672_not ; n15673
g15418 and n15495_not n15672_not ; n15674
g15419 and n15673_not n15674_not ; n15675
g15420 and n15230_not n15234_not ; n15676
g15421 and b[38] n3638 ; n15677
g15422 and b[36] n3843 ; n15678
g15423 and b[37] n3633 ; n15679
g15424 and n15678_not n15679_not ; n15680
g15425 and n15677_not n15680 ; n15681
g15426 and n3641_not n15681 ; n15682
g15427 and n5205_not n15681 ; n15683
g15428 and n15682_not n15683_not ; n15684
g15429 and a[32] n15684_not ; n15685
g15430 and a[32]_not n15684 ; n15686
g15431 and n15685_not n15686_not ; n15687
g15432 and n15676_not n15687_not ; n15688
g15433 and n15676 n15687 ; n15689
g15434 and n15688_not n15689_not ; n15690
g15435 and n15675_not n15690 ; n15691
g15436 and n15675_not n15691_not ; n15692
g15437 and n15690 n15691_not ; n15693
g15438 and n15692_not n15693_not ; n15694
g15439 and n15484 n15694_not ; n15695
g15440 and n15484 n15695_not ; n15696
g15441 and n15694_not n15695_not ; n15697
g15442 and n15696_not n15697_not ; n15698
g15443 and n15253_not n15257_not ; n15699
g15444 and b[44] n2539 ; n15700
g15445 and b[42] n2685 ; n15701
g15446 and b[43] n2534 ; n15702
g15447 and n15701_not n15702_not ; n15703
g15448 and n15700_not n15703 ; n15704
g15449 and n2542_not n15704 ; n15705
g15450 and n7072_not n15704 ; n15706
g15451 and n15705_not n15706_not ; n15707
g15452 and a[26] n15707_not ; n15708
g15453 and a[26]_not n15707 ; n15709
g15454 and n15708_not n15709_not ; n15710
g15455 and n15699_not n15710_not ; n15711
g15456 and n15699_not n15711_not ; n15712
g15457 and n15710_not n15711_not ; n15713
g15458 and n15712_not n15713_not ; n15714
g15459 and n15698_not n15714_not ; n15715
g15460 and n15698_not n15715_not ; n15716
g15461 and n15714_not n15715_not ; n15717
g15462 and n15716_not n15717_not ; n15718
g15463 and n15469 n15718_not ; n15719
g15464 and n15469 n15719_not ; n15720
g15465 and n15718_not n15719_not ; n15721
g15466 and n15720_not n15721_not ; n15722
g15467 and n15454_not n15722 ; n15723
g15468 and n15454 n15722_not ; n15724
g15469 and n15723_not n15724_not ; n15725
g15470 and n15437 n15725_not ; n15726
g15471 and n15437 n15726_not ; n15727
g15472 and n15725_not n15726_not ; n15728
g15473 and n15727_not n15728_not ; n15729
g15474 and n15422_not n15729 ; n15730
g15475 and n15422 n15729_not ; n15731
g15476 and n15730_not n15731_not ; n15732
g15477 and n15405 n15732_not ; n15733
g15478 and n15405 n15733_not ; n15734
g15479 and n15732_not n15733_not ; n15735
g15480 and n15734_not n15735_not ; n15736
g15481 and n15323_not n15327_not ; n15737
g15482 and b[62] n511 ; n15738
g15483 and b[60] n541 ; n15739
g15484 and b[61] n506 ; n15740
g15485 and n15739_not n15740_not ; n15741
g15486 and n15738_not n15741 ; n15742
g15487 and n514_not n15742 ; n15743
g15488 and n13370_not n15742 ; n15744
g15489 and n15743_not n15744_not ; n15745
g15490 and a[8] n15745_not ; n15746
g15491 and a[8]_not n15745 ; n15747
g15492 and n15746_not n15747_not ; n15748
g15493 and n15737_not n15748_not ; n15749
g15494 and n15737_not n15749_not ; n15750
g15495 and n15748_not n15749_not ; n15751
g15496 and n15750_not n15751_not ; n15752
g15497 and n15736_not n15752_not ; n15753
g15498 and n15736 n15751_not ; n15754
g15499 and n15750_not n15754 ; n15755
g15500 and n15753_not n15755_not ; n15756
g15501 and n15390_not n15756 ; n15757
g15502 and n15390 n15756_not ; n15758
g15503 and n15757_not n15758_not ; n15759
g15504 and n15378_not n15759 ; n15760
g15505 and n15378_not n15760_not ; n15761
g15506 and n15759 n15760_not ; n15762
g15507 and n15761_not n15762_not ; n15763
g15508 and n15377_not n15763_not ; n15764
g15509 and n15377 n15762_not ; n15765
g15510 and n15761_not n15765 ; n15766
g15511 and n15764_not n15766_not ; f[68]
g15512 and n15760_not n15764_not ; n15768
g15513 and n15387_not n15757_not ; n15769
g15514 and n15749_not n15753_not ; n15770
g15515 and b[63] n511 ; n15771
g15516 and b[61] n541 ; n15772
g15517 and b[62] n506 ; n15773
g15518 and n15772_not n15773_not ; n15774
g15519 and n15771_not n15774 ; n15775
g15520 and n514 n13771 ; n15776
g15521 and n15775 n15776_not ; n15777
g15522 and a[8] n15777_not ; n15778
g15523 and a[8] n15778_not ; n15779
g15524 and n15777_not n15778_not ; n15780
g15525 and n15779_not n15780_not ; n15781
g15526 and n15770_not n15781_not ; n15782
g15527 and n15770_not n15782_not ; n15783
g15528 and n15781_not n15782_not ; n15784
g15529 and n15783_not n15784_not ; n15785
g15530 and b[60] n700 ; n15786
g15531 and b[58] n767 ; n15787
g15532 and b[59] n695 ; n15788
g15533 and n15787_not n15788_not ; n15789
g15534 and n15786_not n15789 ; n15790
g15535 and n703 n12211 ; n15791
g15536 and n15790 n15791_not ; n15792
g15537 and a[11] n15792_not ; n15793
g15538 and a[11] n15793_not ; n15794
g15539 and n15792_not n15793_not ; n15795
g15540 and n15794_not n15795_not ; n15796
g15541 and n15404_not n15733_not ; n15797
g15542 and n15796 n15797 ; n15798
g15543 and n15796_not n15797_not ; n15799
g15544 and n15798_not n15799_not ; n15800
g15545 and n15435_not n15726_not ; n15801
g15546 and b[54] n1302 ; n15802
g15547 and b[52] n1391 ; n15803
g15548 and b[53] n1297 ; n15804
g15549 and n15803_not n15804_not ; n15805
g15550 and n15802_not n15805 ; n15806
g15551 and n1305 n9998 ; n15807
g15552 and n15806 n15807_not ; n15808
g15553 and a[17] n15808_not ; n15809
g15554 and a[17] n15809_not ; n15810
g15555 and n15808_not n15809_not ; n15811
g15556 and n15810_not n15811_not ; n15812
g15557 and n15801_not n15812_not ; n15813
g15558 and n15801_not n15813_not ; n15814
g15559 and n15812_not n15813_not ; n15815
g15560 and n15814_not n15815_not ; n15816
g15561 and b[48] n2048 ; n15817
g15562 and b[46] n2198 ; n15818
g15563 and b[47] n2043 ; n15819
g15564 and n15818_not n15819_not ; n15820
g15565 and n15817_not n15820 ; n15821
g15566 and n2051 n8009 ; n15822
g15567 and n15821 n15822_not ; n15823
g15568 and a[23] n15823_not ; n15824
g15569 and a[23] n15824_not ; n15825
g15570 and n15823_not n15824_not ; n15826
g15571 and n15825_not n15826_not ; n15827
g15572 and n15468_not n15719_not ; n15828
g15573 and n15827 n15828 ; n15829
g15574 and n15827_not n15828_not ; n15830
g15575 and n15829_not n15830_not ; n15831
g15576 and n15711_not n15715_not ; n15832
g15577 and b[45] n2539 ; n15833
g15578 and b[43] n2685 ; n15834
g15579 and b[44] n2534 ; n15835
g15580 and n15834_not n15835_not ; n15836
g15581 and n15833_not n15836 ; n15837
g15582 and n2542 n7361 ; n15838
g15583 and n15837 n15838_not ; n15839
g15584 and a[26] n15839_not ; n15840
g15585 and a[26] n15840_not ; n15841
g15586 and n15839_not n15840_not ; n15842
g15587 and n15841_not n15842_not ; n15843
g15588 and n15832_not n15843_not ; n15844
g15589 and n15832_not n15844_not ; n15845
g15590 and n15843_not n15844_not ; n15846
g15591 and n15845_not n15846_not ; n15847
g15592 and b[42] n3050 ; n15848
g15593 and b[40] n3243 ; n15849
g15594 and b[41] n3045 ; n15850
g15595 and n15849_not n15850_not ; n15851
g15596 and n15848_not n15851 ; n15852
g15597 and n3053 n6489 ; n15853
g15598 and n15852 n15853_not ; n15854
g15599 and a[29] n15854_not ; n15855
g15600 and a[29] n15855_not ; n15856
g15601 and n15854_not n15855_not ; n15857
g15602 and n15856_not n15857_not ; n15858
g15603 and n15483_not n15695_not ; n15859
g15604 and n15858 n15859 ; n15860
g15605 and n15858_not n15859_not ; n15861
g15606 and n15860_not n15861_not ; n15862
g15607 and n15669_not n15672_not ; n15863
g15608 and n15652_not n15666_not ; n15864
g15609 and n15633_not n15646_not ; n15865
g15610 and n15605_not n15608_not ; n15866
g15611 and n15588_not n15602_not ; n15867
g15612 and n15542_not n15556_not ; n15868
g15613 and b[12] n11531 ; n15869
g15614 and b[10] n11896 ; n15870
g15615 and b[11] n11526 ; n15871
g15616 and n15870_not n15871_not ; n15872
g15617 and n15869_not n15872 ; n15873
g15618 and n842 n11534 ; n15874
g15619 and n15873 n15874_not ; n15875
g15620 and a[59] n15875_not ; n15876
g15621 and a[59] n15876_not ; n15877
g15622 and n15875_not n15876_not ; n15878
g15623 and n15877_not n15878_not ; n15879
g15624 and n15532_not n15536_not ; n15880
g15625 and b[5] n13903 ; n15881
g15626 and b[6] n13488_not ; n15882
g15627 and n15881_not n15882_not ; n15883
g15628 and a[2] a[5]_not ; n15884
g15629 and a[2]_not a[5] ; n15885
g15630 and n15884_not n15885_not ; n15886
g15631 and n15883_not n15886_not ; n15887
g15632 and n15883 n15886 ; n15888
g15633 and n15887_not n15888_not ; n15889
g15634 and n15880 n15889_not ; n15890
g15635 and n15880_not n15889 ; n15891
g15636 and n15890_not n15891_not ; n15892
g15637 and b[9] n12668 ; n15893
g15638 and b[7] n13047 ; n15894
g15639 and b[8] n12663 ; n15895
g15640 and n15894_not n15895_not ; n15896
g15641 and n15893_not n15896 ; n15897
g15642 and n651 n12671 ; n15898
g15643 and n15897 n15898_not ; n15899
g15644 and a[62] n15899_not ; n15900
g15645 and a[62] n15900_not ; n15901
g15646 and n15899_not n15900_not ; n15902
g15647 and n15901_not n15902_not ; n15903
g15648 and n15892_not n15903 ; n15904
g15649 and n15892 n15903_not ; n15905
g15650 and n15904_not n15905_not ; n15906
g15651 and n15879_not n15906 ; n15907
g15652 and n15879_not n15907_not ; n15908
g15653 and n15906 n15907_not ; n15909
g15654 and n15908_not n15909_not ; n15910
g15655 and n15868_not n15910_not ; n15911
g15656 and n15868_not n15911_not ; n15912
g15657 and n15910_not n15911_not ; n15913
g15658 and n15912_not n15913_not ; n15914
g15659 and b[15] n10426 ; n15915
g15660 and b[13] n10796 ; n15916
g15661 and b[14] n10421 ; n15917
g15662 and n15916_not n15917_not ; n15918
g15663 and n15915_not n15918 ; n15919
g15664 and n1131 n10429 ; n15920
g15665 and n15919 n15920_not ; n15921
g15666 and a[56] n15921_not ; n15922
g15667 and a[56] n15922_not ; n15923
g15668 and n15921_not n15922_not ; n15924
g15669 and n15923_not n15924_not ; n15925
g15670 and n15914_not n15925_not ; n15926
g15671 and n15914_not n15926_not ; n15927
g15672 and n15925_not n15926_not ; n15928
g15673 and n15927_not n15928_not ; n15929
g15674 and n15559_not n15562_not ; n15930
g15675 and n15929 n15930 ; n15931
g15676 and n15929_not n15930_not ; n15932
g15677 and n15931_not n15932_not ; n15933
g15678 and b[18] n9339 ; n15934
g15679 and b[16] n9732 ; n15935
g15680 and b[17] n9334 ; n15936
g15681 and n15935_not n15936_not ; n15937
g15682 and n15934_not n15937 ; n15938
g15683 and n1566 n9342 ; n15939
g15684 and n15938 n15939_not ; n15940
g15685 and a[53] n15940_not ; n15941
g15686 and a[53] n15941_not ; n15942
g15687 and n15940_not n15941_not ; n15943
g15688 and n15942_not n15943_not ; n15944
g15689 and n15933 n15944_not ; n15945
g15690 and n15933 n15945_not ; n15946
g15691 and n15944_not n15945_not ; n15947
g15692 and n15946_not n15947_not ; n15948
g15693 and n15567_not n15582_not ; n15949
g15694 and n15948 n15949 ; n15950
g15695 and n15948_not n15949_not ; n15951
g15696 and n15950_not n15951_not ; n15952
g15697 and b[21] n8362 ; n15953
g15698 and b[19] n8715 ; n15954
g15699 and b[20] n8357 ; n15955
g15700 and n15954_not n15955_not ; n15956
g15701 and n15953_not n15956 ; n15957
g15702 and n1984 n8365 ; n15958
g15703 and n15957 n15958_not ; n15959
g15704 and a[50] n15959_not ; n15960
g15705 and a[50] n15960_not ; n15961
g15706 and n15959_not n15960_not ; n15962
g15707 and n15961_not n15962_not ; n15963
g15708 and n15952 n15963_not ; n15964
g15709 and n15952 n15964_not ; n15965
g15710 and n15963_not n15964_not ; n15966
g15711 and n15965_not n15966_not ; n15967
g15712 and n15867_not n15967 ; n15968
g15713 and n15867 n15967_not ; n15969
g15714 and n15968_not n15969_not ; n15970
g15715 and b[24] n7446 ; n15971
g15716 and b[22] n7787 ; n15972
g15717 and b[23] n7441 ; n15973
g15718 and n15972_not n15973_not ; n15974
g15719 and n15971_not n15974 ; n15975
g15720 and n2458 n7449 ; n15976
g15721 and n15975 n15976_not ; n15977
g15722 and a[47] n15977_not ; n15978
g15723 and a[47] n15978_not ; n15979
g15724 and n15977_not n15978_not ; n15980
g15725 and n15979_not n15980_not ; n15981
g15726 and n15970_not n15981_not ; n15982
g15727 and n15970 n15981 ; n15983
g15728 and n15982_not n15983_not ; n15984
g15729 and n15866 n15984_not ; n15985
g15730 and n15866_not n15984 ; n15986
g15731 and n15985_not n15986_not ; n15987
g15732 and b[27] n6595 ; n15988
g15733 and b[25] n6902 ; n15989
g15734 and b[26] n6590 ; n15990
g15735 and n15989_not n15990_not ; n15991
g15736 and n15988_not n15991 ; n15992
g15737 and n2990 n6598 ; n15993
g15738 and n15992 n15993_not ; n15994
g15739 and a[44] n15994_not ; n15995
g15740 and a[44] n15995_not ; n15996
g15741 and n15994_not n15995_not ; n15997
g15742 and n15996_not n15997_not ; n15998
g15743 and n15987 n15998_not ; n15999
g15744 and n15987 n15999_not ; n16000
g15745 and n15998_not n15999_not ; n16001
g15746 and n16000_not n16001_not ; n16002
g15747 and n15614_not n15627_not ; n16003
g15748 and n16002 n16003 ; n16004
g15749 and n16002_not n16003_not ; n16005
g15750 and n16004_not n16005_not ; n16006
g15751 and b[30] n5777 ; n16007
g15752 and b[28] n6059 ; n16008
g15753 and b[29] n5772 ; n16009
g15754 and n16008_not n16009_not ; n16010
g15755 and n16007_not n16010 ; n16011
g15756 and n3577 n5780 ; n16012
g15757 and n16011 n16012_not ; n16013
g15758 and a[41] n16013_not ; n16014
g15759 and a[41] n16014_not ; n16015
g15760 and n16013_not n16014_not ; n16016
g15761 and n16015_not n16016_not ; n16017
g15762 and n16006 n16017_not ; n16018
g15763 and n16006_not n16017 ; n16019
g15764 and n15865_not n16019_not ; n16020
g15765 and n16018_not n16020 ; n16021
g15766 and n15865_not n16021_not ; n16022
g15767 and n16018_not n16021_not ; n16023
g15768 and n16019_not n16023 ; n16024
g15769 and n16022_not n16024_not ; n16025
g15770 and b[33] n5035 ; n16026
g15771 and b[31] n5277 ; n16027
g15772 and b[32] n5030 ; n16028
g15773 and n16027_not n16028_not ; n16029
g15774 and n16026_not n16029 ; n16030
g15775 and n4223 n5038 ; n16031
g15776 and n16030 n16031_not ; n16032
g15777 and a[38] n16032_not ; n16033
g15778 and a[38] n16033_not ; n16034
g15779 and n16032_not n16033_not ; n16035
g15780 and n16034_not n16035_not ; n16036
g15781 and n16025_not n16036_not ; n16037
g15782 and n16025_not n16037_not ; n16038
g15783 and n16036_not n16037_not ; n16039
g15784 and n16038_not n16039_not ; n16040
g15785 and n15864_not n16040 ; n16041
g15786 and n15864 n16040_not ; n16042
g15787 and n16041_not n16042_not ; n16043
g15788 and b[36] n4287 ; n16044
g15789 and b[34] n4532 ; n16045
g15790 and b[35] n4282 ; n16046
g15791 and n16045_not n16046_not ; n16047
g15792 and n16044_not n16047 ; n16048
g15793 and n4290 n4922 ; n16049
g15794 and n16048 n16049_not ; n16050
g15795 and a[35] n16050_not ; n16051
g15796 and a[35] n16051_not ; n16052
g15797 and n16050_not n16051_not ; n16053
g15798 and n16052_not n16053_not ; n16054
g15799 and n16043_not n16054_not ; n16055
g15800 and n16043 n16054 ; n16056
g15801 and n16055_not n16056_not ; n16057
g15802 and n15863 n16057_not ; n16058
g15803 and n15863_not n16057 ; n16059
g15804 and n16058_not n16059_not ; n16060
g15805 and b[39] n3638 ; n16061
g15806 and b[37] n3843 ; n16062
g15807 and b[38] n3633 ; n16063
g15808 and n16062_not n16063_not ; n16064
g15809 and n16061_not n16064 ; n16065
g15810 and n3641 n5451 ; n16066
g15811 and n16065 n16066_not ; n16067
g15812 and a[32] n16067_not ; n16068
g15813 and a[32] n16068_not ; n16069
g15814 and n16067_not n16068_not ; n16070
g15815 and n16069_not n16070_not ; n16071
g15816 and n15688_not n15691_not ; n16072
g15817 and n16071 n16072 ; n16073
g15818 and n16071_not n16072_not ; n16074
g15819 and n16073_not n16074_not ; n16075
g15820 and n16060 n16075 ; n16076
g15821 and n16060_not n16075_not ; n16077
g15822 and n16076_not n16077_not ; n16078
g15823 and n15862 n16078 ; n16079
g15824 and n15862_not n16078_not ; n16080
g15825 and n16079_not n16080_not ; n16081
g15826 and n15847_not n16081_not ; n16082
g15827 and n15847 n16081 ; n16083
g15828 and n16082_not n16083_not ; n16084
g15829 and n15831 n16084_not ; n16085
g15830 and n15831 n16085_not ; n16086
g15831 and n16084_not n16085_not ; n16087
g15832 and n16086_not n16087_not ; n16088
g15833 and b[51] n1627 ; n16089
g15834 and b[49] n1763 ; n16090
g15835 and b[50] n1622 ; n16091
g15836 and n16090_not n16091_not ; n16092
g15837 and n16089_not n16092 ; n16093
g15838 and n1630 n8976 ; n16094
g15839 and n16093 n16094_not ; n16095
g15840 and a[20] n16095_not ; n16096
g15841 and a[20] n16096_not ; n16097
g15842 and n16095_not n16096_not ; n16098
g15843 and n16097_not n16098_not ; n16099
g15844 and n15454_not n15722_not ; n16100
g15845 and n15451_not n16100_not ; n16101
g15846 and n16099_not n16101_not ; n16102
g15847 and n16099 n16101 ; n16103
g15848 and n16102_not n16103_not ; n16104
g15849 and n16088_not n16104 ; n16105
g15850 and n16088_not n16105_not ; n16106
g15851 and n16104 n16105_not ; n16107
g15852 and n16106_not n16107_not ; n16108
g15853 and n15816_not n16108_not ; n16109
g15854 and n15816_not n16109_not ; n16110
g15855 and n16108_not n16109_not ; n16111
g15856 and n16110_not n16111_not ; n16112
g15857 and b[57] n951 ; n16113
g15858 and b[55] n1056 ; n16114
g15859 and b[56] n946 ; n16115
g15860 and n16114_not n16115_not ; n16116
g15861 and n16113_not n16116 ; n16117
g15862 and n954 n11410 ; n16118
g15863 and n16117 n16118_not ; n16119
g15864 and a[14] n16119_not ; n16120
g15865 and a[14] n16120_not ; n16121
g15866 and n16119_not n16120_not ; n16122
g15867 and n16121_not n16122_not ; n16123
g15868 and n15422_not n15729_not ; n16124
g15869 and n15419_not n16124_not ; n16125
g15870 and n16123_not n16125_not ; n16126
g15871 and n16123 n16125 ; n16127
g15872 and n16126_not n16127_not ; n16128
g15873 and n16112_not n16128 ; n16129
g15874 and n16112_not n16129_not ; n16130
g15875 and n16128 n16129_not ; n16131
g15876 and n16130_not n16131_not ; n16132
g15877 and n15800 n16132_not ; n16133
g15878 and n15800 n16133_not ; n16134
g15879 and n16132_not n16133_not ; n16135
g15880 and n16134_not n16135_not ; n16136
g15881 and n15785_not n16136 ; n16137
g15882 and n15785 n16136_not ; n16138
g15883 and n16137_not n16138_not ; n16139
g15884 and n15769_not n16139_not ; n16140
g15885 and n15769 n16139 ; n16141
g15886 and n16140_not n16141_not ; n16142
g15887 and n15768_not n16142 ; n16143
g15888 and n15768 n16142_not ; n16144
g15889 and n16143_not n16144_not ; f[69]
g15890 and n15799_not n16133_not ; n16146
g15891 and b[62] n541 ; n16147
g15892 and b[63] n506 ; n16148
g15893 and n16147_not n16148_not ; n16149
g15894 and n514_not n16149 ; n16150
g15895 and n13800 n16149 ; n16151
g15896 and n16150_not n16151_not ; n16152
g15897 and a[8] n16152_not ; n16153
g15898 and a[8]_not n16152 ; n16154
g15899 and n16153_not n16154_not ; n16155
g15900 and n16146_not n16155_not ; n16156
g15901 and n16146 n16155 ; n16157
g15902 and n16156_not n16157_not ; n16158
g15903 and b[61] n700 ; n16159
g15904 and b[59] n767 ; n16160
g15905 and b[60] n695 ; n16161
g15906 and n16160_not n16161_not ; n16162
g15907 and n16159_not n16162 ; n16163
g15908 and n703 n12969 ; n16164
g15909 and n16163 n16164_not ; n16165
g15910 and a[11] n16165_not ; n16166
g15911 and a[11] n16166_not ; n16167
g15912 and n16165_not n16166_not ; n16168
g15913 and n16167_not n16168_not ; n16169
g15914 and n16126_not n16129_not ; n16170
g15915 and n16169 n16170 ; n16171
g15916 and n16169_not n16170_not ; n16172
g15917 and n16171_not n16172_not ; n16173
g15918 and n15813_not n16109_not ; n16174
g15919 and b[58] n951 ; n16175
g15920 and b[56] n1056 ; n16176
g15921 and b[57] n946 ; n16177
g15922 and n16176_not n16177_not ; n16178
g15923 and n16175_not n16178 ; n16179
g15924 and n954_not n16179 ; n16180
g15925 and n11436_not n16179 ; n16181
g15926 and n16180_not n16181_not ; n16182
g15927 and a[14] n16182_not ; n16183
g15928 and a[14]_not n16182 ; n16184
g15929 and n16183_not n16184_not ; n16185
g15930 and n16174_not n16185_not ; n16186
g15931 and n16174 n16185 ; n16187
g15932 and n16186_not n16187_not ; n16188
g15933 and b[55] n1302 ; n16189
g15934 and b[53] n1391 ; n16190
g15935 and b[54] n1297 ; n16191
g15936 and n16190_not n16191_not ; n16192
g15937 and n16189_not n16192 ; n16193
g15938 and n1305 n10684 ; n16194
g15939 and n16193 n16194_not ; n16195
g15940 and a[17] n16195_not ; n16196
g15941 and a[17] n16196_not ; n16197
g15942 and n16195_not n16196_not ; n16198
g15943 and n16197_not n16198_not ; n16199
g15944 and n16102_not n16105_not ; n16200
g15945 and n16199 n16200 ; n16201
g15946 and n16199_not n16200_not ; n16202
g15947 and n16201_not n16202_not ; n16203
g15948 and b[52] n1627 ; n16204
g15949 and b[50] n1763 ; n16205
g15950 and b[51] n1622 ; n16206
g15951 and n16205_not n16206_not ; n16207
g15952 and n16204_not n16207 ; n16208
g15953 and n1630 n9628 ; n16209
g15954 and n16208 n16209_not ; n16210
g15955 and a[20] n16210_not ; n16211
g15956 and a[20] n16211_not ; n16212
g15957 and n16210_not n16211_not ; n16213
g15958 and n16212_not n16213_not ; n16214
g15959 and n15830_not n16085_not ; n16215
g15960 and n16214 n16215 ; n16216
g15961 and n16214_not n16215_not ; n16217
g15962 and n16216_not n16217_not ; n16218
g15963 and b[49] n2048 ; n16219
g15964 and b[47] n2198 ; n16220
g15965 and b[48] n2043 ; n16221
g15966 and n16220_not n16221_not ; n16222
g15967 and n16219_not n16222 ; n16223
g15968 and n2051 n8625 ; n16224
g15969 and n16223 n16224_not ; n16225
g15970 and a[23] n16225_not ; n16226
g15971 and a[23] n16226_not ; n16227
g15972 and n16225_not n16226_not ; n16228
g15973 and n16227_not n16228_not ; n16229
g15974 and n15847_not n16081 ; n16230
g15975 and n15844_not n16230_not ; n16231
g15976 and n16229_not n16231_not ; n16232
g15977 and n16229_not n16232_not ; n16233
g15978 and n16231_not n16232_not ; n16234
g15979 and n16233_not n16234_not ; n16235
g15980 and n15861_not n16079_not ; n16236
g15981 and b[46] n2539 ; n16237
g15982 and b[44] n2685 ; n16238
g15983 and b[45] n2534 ; n16239
g15984 and n16238_not n16239_not ; n16240
g15985 and n16237_not n16240 ; n16241
g15986 and n2542_not n16241 ; n16242
g15987 and n7677_not n16241 ; n16243
g15988 and n16242_not n16243_not ; n16244
g15989 and a[26] n16244_not ; n16245
g15990 and a[26]_not n16244 ; n16246
g15991 and n16245_not n16246_not ; n16247
g15992 and n16236_not n16247_not ; n16248
g15993 and n16236 n16247 ; n16249
g15994 and n16248_not n16249_not ; n16250
g15995 and b[43] n3050 ; n16251
g15996 and b[41] n3243 ; n16252
g15997 and b[42] n3045 ; n16253
g15998 and n16252_not n16253_not ; n16254
g15999 and n16251_not n16254 ; n16255
g16000 and n3053 n6515 ; n16256
g16001 and n16255 n16256_not ; n16257
g16002 and a[29] n16257_not ; n16258
g16003 and a[29] n16258_not ; n16259
g16004 and n16257_not n16258_not ; n16260
g16005 and n16259_not n16260_not ; n16261
g16006 and n16074_not n16076_not ; n16262
g16007 and n16261_not n16262_not ; n16263
g16008 and n16261_not n16263_not ; n16264
g16009 and n16262_not n16263_not ; n16265
g16010 and n16264_not n16265_not ; n16266
g16011 and b[40] n3638 ; n16267
g16012 and b[38] n3843 ; n16268
g16013 and b[39] n3633 ; n16269
g16014 and n16268_not n16269_not ; n16270
g16015 and n16267_not n16270 ; n16271
g16016 and n3641 n5955 ; n16272
g16017 and n16271 n16272_not ; n16273
g16018 and a[32] n16273_not ; n16274
g16019 and a[32] n16274_not ; n16275
g16020 and n16273_not n16274_not ; n16276
g16021 and n16275_not n16276_not ; n16277
g16022 and n16055_not n16059_not ; n16278
g16023 and n16277 n16278 ; n16279
g16024 and n16277_not n16278_not ; n16280
g16025 and n16279_not n16280_not ; n16281
g16026 and b[37] n4287 ; n16282
g16027 and b[35] n4532 ; n16283
g16028 and b[36] n4282 ; n16284
g16029 and n16283_not n16284_not ; n16285
g16030 and n16282_not n16285 ; n16286
g16031 and n4290 n5181 ; n16287
g16032 and n16286 n16287_not ; n16288
g16033 and a[35] n16288_not ; n16289
g16034 and a[35] n16289_not ; n16290
g16035 and n16288_not n16289_not ; n16291
g16036 and n16290_not n16291_not ; n16292
g16037 and n15864_not n16040_not ; n16293
g16038 and n16037_not n16293_not ; n16294
g16039 and b[34] n5035 ; n16295
g16040 and b[32] n5277 ; n16296
g16041 and b[33] n5030 ; n16297
g16042 and n16296_not n16297_not ; n16298
g16043 and n16295_not n16298 ; n16299
g16044 and n4466 n5038 ; n16300
g16045 and n16299 n16300_not ; n16301
g16046 and a[38] n16301_not ; n16302
g16047 and a[38] n16302_not ; n16303
g16048 and n16301_not n16302_not ; n16304
g16049 and n16303_not n16304_not ; n16305
g16050 and n15891_not n15905_not ; n16306
g16051 and a[2]_not a[5]_not ; n16307
g16052 and n15887_not n16307_not ; n16308
g16053 and b[6] n13903 ; n16309
g16054 and b[7] n13488_not ; n16310
g16055 and n16309_not n16310_not ; n16311
g16056 and n16308_not n16311 ; n16312
g16057 and n16308 n16311_not ; n16313
g16058 and n16312_not n16313_not ; n16314
g16059 and b[10] n12668 ; n16315
g16060 and b[8] n13047 ; n16316
g16061 and b[9] n12663 ; n16317
g16062 and n16316_not n16317_not ; n16318
g16063 and n16315_not n16318 ; n16319
g16064 and n12671_not n16319 ; n16320
g16065 and n738_not n16319 ; n16321
g16066 and n16320_not n16321_not ; n16322
g16067 and a[62] n16322_not ; n16323
g16068 and a[62]_not n16322 ; n16324
g16069 and n16323_not n16324_not ; n16325
g16070 and n16314 n16325_not ; n16326
g16071 and n16314_not n16325 ; n16327
g16072 and n16326_not n16327_not ; n16328
g16073 and n16306_not n16328 ; n16329
g16074 and n16306 n16328_not ; n16330
g16075 and n16329_not n16330_not ; n16331
g16076 and b[13] n11531 ; n16332
g16077 and b[11] n11896 ; n16333
g16078 and b[12] n11526 ; n16334
g16079 and n16333_not n16334_not ; n16335
g16080 and n16332_not n16335 ; n16336
g16081 and n1008 n11534 ; n16337
g16082 and n16336 n16337_not ; n16338
g16083 and a[59] n16338_not ; n16339
g16084 and a[59] n16339_not ; n16340
g16085 and n16338_not n16339_not ; n16341
g16086 and n16340_not n16341_not ; n16342
g16087 and n16331 n16342_not ; n16343
g16088 and n16331 n16343_not ; n16344
g16089 and n16342_not n16343_not ; n16345
g16090 and n16344_not n16345_not ; n16346
g16091 and n15907_not n15911_not ; n16347
g16092 and n16346 n16347 ; n16348
g16093 and n16346_not n16347_not ; n16349
g16094 and n16348_not n16349_not ; n16350
g16095 and b[16] n10426 ; n16351
g16096 and b[14] n10796 ; n16352
g16097 and b[15] n10421 ; n16353
g16098 and n16352_not n16353_not ; n16354
g16099 and n16351_not n16354 ; n16355
g16100 and n1237 n10429 ; n16356
g16101 and n16355 n16356_not ; n16357
g16102 and a[56] n16357_not ; n16358
g16103 and a[56] n16358_not ; n16359
g16104 and n16357_not n16358_not ; n16360
g16105 and n16359_not n16360_not ; n16361
g16106 and n16350 n16361_not ; n16362
g16107 and n16350 n16362_not ; n16363
g16108 and n16361_not n16362_not ; n16364
g16109 and n16363_not n16364_not ; n16365
g16110 and n15926_not n15932_not ; n16366
g16111 and n16365 n16366 ; n16367
g16112 and n16365_not n16366_not ; n16368
g16113 and n16367_not n16368_not ; n16369
g16114 and b[19] n9339 ; n16370
g16115 and b[17] n9732 ; n16371
g16116 and b[18] n9334 ; n16372
g16117 and n16371_not n16372_not ; n16373
g16118 and n16370_not n16373 ; n16374
g16119 and n1708 n9342 ; n16375
g16120 and n16374 n16375_not ; n16376
g16121 and a[53] n16376_not ; n16377
g16122 and a[53] n16377_not ; n16378
g16123 and n16376_not n16377_not ; n16379
g16124 and n16378_not n16379_not ; n16380
g16125 and n16369 n16380_not ; n16381
g16126 and n16369 n16381_not ; n16382
g16127 and n16380_not n16381_not ; n16383
g16128 and n16382_not n16383_not ; n16384
g16129 and n15945_not n15951_not ; n16385
g16130 and n16384 n16385 ; n16386
g16131 and n16384_not n16385_not ; n16387
g16132 and n16386_not n16387_not ; n16388
g16133 and b[22] n8362 ; n16389
g16134 and b[20] n8715 ; n16390
g16135 and b[21] n8357 ; n16391
g16136 and n16390_not n16391_not ; n16392
g16137 and n16389_not n16392 ; n16393
g16138 and n2145 n8365 ; n16394
g16139 and n16393 n16394_not ; n16395
g16140 and a[50] n16395_not ; n16396
g16141 and a[50] n16396_not ; n16397
g16142 and n16395_not n16396_not ; n16398
g16143 and n16397_not n16398_not ; n16399
g16144 and n16388 n16399_not ; n16400
g16145 and n16388 n16400_not ; n16401
g16146 and n16399_not n16400_not ; n16402
g16147 and n16401_not n16402_not ; n16403
g16148 and n15867_not n15967_not ; n16404
g16149 and n15964_not n16404_not ; n16405
g16150 and n16403 n16405 ; n16406
g16151 and n16403_not n16405_not ; n16407
g16152 and n16406_not n16407_not ; n16408
g16153 and b[25] n7446 ; n16409
g16154 and b[23] n7787 ; n16410
g16155 and b[24] n7441 ; n16411
g16156 and n16410_not n16411_not ; n16412
g16157 and n16409_not n16412 ; n16413
g16158 and n2485 n7449 ; n16414
g16159 and n16413 n16414_not ; n16415
g16160 and a[47] n16415_not ; n16416
g16161 and a[47] n16416_not ; n16417
g16162 and n16415_not n16416_not ; n16418
g16163 and n16417_not n16418_not ; n16419
g16164 and n16408 n16419_not ; n16420
g16165 and n16408 n16420_not ; n16421
g16166 and n16419_not n16420_not ; n16422
g16167 and n16421_not n16422_not ; n16423
g16168 and n15982_not n15986_not ; n16424
g16169 and n16423 n16424 ; n16425
g16170 and n16423_not n16424_not ; n16426
g16171 and n16425_not n16426_not ; n16427
g16172 and b[28] n6595 ; n16428
g16173 and b[26] n6902 ; n16429
g16174 and b[27] n6590 ; n16430
g16175 and n16429_not n16430_not ; n16431
g16176 and n16428_not n16431 ; n16432
g16177 and n3189 n6598 ; n16433
g16178 and n16432 n16433_not ; n16434
g16179 and a[44] n16434_not ; n16435
g16180 and a[44] n16435_not ; n16436
g16181 and n16434_not n16435_not ; n16437
g16182 and n16436_not n16437_not ; n16438
g16183 and n16427 n16438_not ; n16439
g16184 and n16427 n16439_not ; n16440
g16185 and n16438_not n16439_not ; n16441
g16186 and n16440_not n16441_not ; n16442
g16187 and n15999_not n16005_not ; n16443
g16188 and n16442 n16443 ; n16444
g16189 and n16442_not n16443_not ; n16445
g16190 and n16444_not n16445_not ; n16446
g16191 and b[31] n5777 ; n16447
g16192 and b[29] n6059 ; n16448
g16193 and b[30] n5772 ; n16449
g16194 and n16448_not n16449_not ; n16450
g16195 and n16447_not n16450 ; n16451
g16196 and n3796 n5780 ; n16452
g16197 and n16451 n16452_not ; n16453
g16198 and a[41] n16453_not ; n16454
g16199 and a[41] n16454_not ; n16455
g16200 and n16453_not n16454_not ; n16456
g16201 and n16455_not n16456_not ; n16457
g16202 and n16446_not n16457 ; n16458
g16203 and n16446 n16457_not ; n16459
g16204 and n16458_not n16459_not ; n16460
g16205 and n16023_not n16460 ; n16461
g16206 and n16023 n16460_not ; n16462
g16207 and n16461_not n16462_not ; n16463
g16208 and n16305_not n16463 ; n16464
g16209 and n16305 n16463_not ; n16465
g16210 and n16464_not n16465_not ; n16466
g16211 and n16294_not n16466 ; n16467
g16212 and n16294 n16466_not ; n16468
g16213 and n16467_not n16468_not ; n16469
g16214 and n16292_not n16469 ; n16470
g16215 and n16292_not n16470_not ; n16471
g16216 and n16469 n16470_not ; n16472
g16217 and n16471_not n16472_not ; n16473
g16218 and n16281 n16473_not ; n16474
g16219 and n16281 n16474_not ; n16475
g16220 and n16473_not n16474_not ; n16476
g16221 and n16475_not n16476_not ; n16477
g16222 and n16266_not n16477 ; n16478
g16223 and n16266 n16477_not ; n16479
g16224 and n16478_not n16479_not ; n16480
g16225 and n16250 n16480_not ; n16481
g16226 and n16250 n16481_not ; n16482
g16227 and n16480_not n16481_not ; n16483
g16228 and n16482_not n16483_not ; n16484
g16229 and n16235_not n16484 ; n16485
g16230 and n16235 n16484_not ; n16486
g16231 and n16485_not n16486_not ; n16487
g16232 and n16218 n16487_not ; n16488
g16233 and n16218 n16488_not ; n16489
g16234 and n16487_not n16488_not ; n16490
g16235 and n16489_not n16490_not ; n16491
g16236 and n16203 n16491_not ; n16492
g16237 and n16203_not n16491 ; n16493
g16238 and n16188 n16493_not ; n16494
g16239 and n16492_not n16494 ; n16495
g16240 and n16188 n16495_not ; n16496
g16241 and n16493_not n16495_not ; n16497
g16242 and n16492_not n16497 ; n16498
g16243 and n16496_not n16498_not ; n16499
g16244 and n16173 n16499_not ; n16500
g16245 and n16173_not n16499 ; n16501
g16246 and n16158 n16501_not ; n16502
g16247 and n16500_not n16502 ; n16503
g16248 and n16158 n16503_not ; n16504
g16249 and n16501_not n16503_not ; n16505
g16250 and n16500_not n16505 ; n16506
g16251 and n16504_not n16506_not ; n16507
g16252 and n15785_not n16136_not ; n16508
g16253 and n15782_not n16508_not ; n16509
g16254 and n16507_not n16509_not ; n16510
g16255 and n16507_not n16510_not ; n16511
g16256 and n16509_not n16510_not ; n16512
g16257 and n16511_not n16512_not ; n16513
g16258 and n16140_not n16143_not ; n16514
g16259 and n16513_not n16514_not ; n16515
g16260 and n16513 n16514 ; n16516
g16261 and n16515_not n16516_not ; f[70]
g16262 and n16510_not n16515_not ; n16518
g16263 and n16156_not n16503_not ; n16519
g16264 and n16172_not n16500_not ; n16520
g16265 and b[63] n541 ; n16521
g16266 and n514 n13797 ; n16522
g16267 and n16521_not n16522_not ; n16523
g16268 and a[8] n16523_not ; n16524
g16269 and a[8] n16524_not ; n16525
g16270 and n16523_not n16524_not ; n16526
g16271 and n16525_not n16526_not ; n16527
g16272 and n16520_not n16527_not ; n16528
g16273 and n16520_not n16528_not ; n16529
g16274 and n16527_not n16528_not ; n16530
g16275 and n16529_not n16530_not ; n16531
g16276 and b[56] n1302 ; n16532
g16277 and b[54] n1391 ; n16533
g16278 and b[55] n1297 ; n16534
g16279 and n16533_not n16534_not ; n16535
g16280 and n16532_not n16535 ; n16536
g16281 and n1305 n10708 ; n16537
g16282 and n16536 n16537_not ; n16538
g16283 and a[17] n16538_not ; n16539
g16284 and a[17] n16539_not ; n16540
g16285 and n16538_not n16539_not ; n16541
g16286 and n16540_not n16541_not ; n16542
g16287 and n16217_not n16488_not ; n16543
g16288 and n16542 n16543 ; n16544
g16289 and n16542_not n16543_not ; n16545
g16290 and n16544_not n16545_not ; n16546
g16291 and b[50] n2048 ; n16547
g16292 and b[48] n2198 ; n16548
g16293 and b[49] n2043 ; n16549
g16294 and n16548_not n16549_not ; n16550
g16295 and n16547_not n16550 ; n16551
g16296 and n2051 n8949 ; n16552
g16297 and n16551 n16552_not ; n16553
g16298 and a[23] n16553_not ; n16554
g16299 and a[23] n16554_not ; n16555
g16300 and n16553_not n16554_not ; n16556
g16301 and n16555_not n16556_not ; n16557
g16302 and n16248_not n16481_not ; n16558
g16303 and n16557 n16558 ; n16559
g16304 and n16557_not n16558_not ; n16560
g16305 and n16559_not n16560_not ; n16561
g16306 and b[47] n2539 ; n16562
g16307 and b[45] n2685 ; n16563
g16308 and b[46] n2534 ; n16564
g16309 and n16563_not n16564_not ; n16565
g16310 and n16562_not n16565 ; n16566
g16311 and n2542 n7703 ; n16567
g16312 and n16566 n16567_not ; n16568
g16313 and a[26] n16568_not ; n16569
g16314 and a[26] n16569_not ; n16570
g16315 and n16568_not n16569_not ; n16571
g16316 and n16570_not n16571_not ; n16572
g16317 and n16266_not n16477_not ; n16573
g16318 and n16263_not n16573_not ; n16574
g16319 and n16572_not n16574_not ; n16575
g16320 and n16572_not n16575_not ; n16576
g16321 and n16574_not n16575_not ; n16577
g16322 and n16576_not n16577_not ; n16578
g16323 and b[41] n3638 ; n16579
g16324 and b[39] n3843 ; n16580
g16325 and b[40] n3633 ; n16581
g16326 and n16580_not n16581_not ; n16582
g16327 and n16579_not n16582 ; n16583
g16328 and n3641 n6219 ; n16584
g16329 and n16583 n16584_not ; n16585
g16330 and a[32] n16585_not ; n16586
g16331 and a[32] n16586_not ; n16587
g16332 and n16585_not n16586_not ; n16588
g16333 and n16587_not n16588_not ; n16589
g16334 and n16467_not n16470_not ; n16590
g16335 and n16589 n16590 ; n16591
g16336 and n16589_not n16590_not ; n16592
g16337 and n16591_not n16592_not ; n16593
g16338 and b[35] n5035 ; n16594
g16339 and b[33] n5277 ; n16595
g16340 and b[34] n5030 ; n16596
g16341 and n16595_not n16596_not ; n16597
g16342 and n16594_not n16597 ; n16598
g16343 and n4696 n5038 ; n16599
g16344 and n16598 n16599_not ; n16600
g16345 and a[38] n16600_not ; n16601
g16346 and a[38] n16601_not ; n16602
g16347 and n16600_not n16601_not ; n16603
g16348 and n16602_not n16603_not ; n16604
g16349 and b[26] n7446 ; n16605
g16350 and b[24] n7787 ; n16606
g16351 and b[25] n7441 ; n16607
g16352 and n16606_not n16607_not ; n16608
g16353 and n16605_not n16608 ; n16609
g16354 and n2813 n7449 ; n16610
g16355 and n16609 n16610_not ; n16611
g16356 and a[47] n16611_not ; n16612
g16357 and a[47] n16612_not ; n16613
g16358 and n16611_not n16612_not ; n16614
g16359 and n16613_not n16614_not ; n16615
g16360 and n16387_not n16400_not ; n16616
g16361 and b[23] n8362 ; n16617
g16362 and b[21] n8715 ; n16618
g16363 and b[22] n8357 ; n16619
g16364 and n16618_not n16619_not ; n16620
g16365 and n16617_not n16620 ; n16621
g16366 and n2300 n8365 ; n16622
g16367 and n16621 n16622_not ; n16623
g16368 and a[50] n16623_not ; n16624
g16369 and a[50] n16624_not ; n16625
g16370 and n16623_not n16624_not ; n16626
g16371 and n16625_not n16626_not ; n16627
g16372 and n16368_not n16381_not ; n16628
g16373 and n16329_not n16343_not ; n16629
g16374 and n16312_not n16326_not ; n16630
g16375 and b[7] n13903 ; n16631
g16376 and b[8] n13488_not ; n16632
g16377 and n16631_not n16632_not ; n16633
g16378 and n16311 n16633_not ; n16634
g16379 and n16311_not n16633 ; n16635
g16380 and n16630_not n16635_not ; n16636
g16381 and n16634_not n16636 ; n16637
g16382 and n16630_not n16637_not ; n16638
g16383 and n16635_not n16637_not ; n16639
g16384 and n16634_not n16639 ; n16640
g16385 and n16638_not n16640_not ; n16641
g16386 and b[11] n12668 ; n16642
g16387 and b[9] n13047 ; n16643
g16388 and b[10] n12663 ; n16644
g16389 and n16643_not n16644_not ; n16645
g16390 and n16642_not n16645 ; n16646
g16391 and n818 n12671 ; n16647
g16392 and n16646 n16647_not ; n16648
g16393 and a[62] n16648_not ; n16649
g16394 and a[62] n16649_not ; n16650
g16395 and n16648_not n16649_not ; n16651
g16396 and n16650_not n16651_not ; n16652
g16397 and n16641_not n16652 ; n16653
g16398 and n16641 n16652_not ; n16654
g16399 and n16653_not n16654_not ; n16655
g16400 and b[14] n11531 ; n16656
g16401 and b[12] n11896 ; n16657
g16402 and b[13] n11526 ; n16658
g16403 and n16657_not n16658_not ; n16659
g16404 and n16656_not n16659 ; n16660
g16405 and n1034 n11534 ; n16661
g16406 and n16660 n16661_not ; n16662
g16407 and a[59] n16662_not ; n16663
g16408 and a[59] n16663_not ; n16664
g16409 and n16662_not n16663_not ; n16665
g16410 and n16664_not n16665_not ; n16666
g16411 and n16655_not n16666_not ; n16667
g16412 and n16655 n16666 ; n16668
g16413 and n16667_not n16668_not ; n16669
g16414 and n16629 n16669_not ; n16670
g16415 and n16629_not n16669 ; n16671
g16416 and n16670_not n16671_not ; n16672
g16417 and b[17] n10426 ; n16673
g16418 and b[15] n10796 ; n16674
g16419 and b[16] n10421 ; n16675
g16420 and n16674_not n16675_not ; n16676
g16421 and n16673_not n16676 ; n16677
g16422 and n1356 n10429 ; n16678
g16423 and n16677 n16678_not ; n16679
g16424 and a[56] n16679_not ; n16680
g16425 and a[56] n16680_not ; n16681
g16426 and n16679_not n16680_not ; n16682
g16427 and n16681_not n16682_not ; n16683
g16428 and n16672 n16683_not ; n16684
g16429 and n16672 n16684_not ; n16685
g16430 and n16683_not n16684_not ; n16686
g16431 and n16685_not n16686_not ; n16687
g16432 and n16349_not n16362_not ; n16688
g16433 and n16687 n16688 ; n16689
g16434 and n16687_not n16688_not ; n16690
g16435 and n16689_not n16690_not ; n16691
g16436 and b[20] n9339 ; n16692
g16437 and b[18] n9732 ; n16693
g16438 and b[19] n9334 ; n16694
g16439 and n16693_not n16694_not ; n16695
g16440 and n16692_not n16695 ; n16696
g16441 and n1846 n9342 ; n16697
g16442 and n16696 n16697_not ; n16698
g16443 and a[53] n16698_not ; n16699
g16444 and a[53] n16699_not ; n16700
g16445 and n16698_not n16699_not ; n16701
g16446 and n16700_not n16701_not ; n16702
g16447 and n16691_not n16702 ; n16703
g16448 and n16691 n16702_not ; n16704
g16449 and n16703_not n16704_not ; n16705
g16450 and n16628_not n16705 ; n16706
g16451 and n16628_not n16706_not ; n16707
g16452 and n16705 n16706_not ; n16708
g16453 and n16707_not n16708_not ; n16709
g16454 and n16627_not n16709_not ; n16710
g16455 and n16627 n16708_not ; n16711
g16456 and n16707_not n16711 ; n16712
g16457 and n16710_not n16712_not ; n16713
g16458 and n16616_not n16713 ; n16714
g16459 and n16616 n16713_not ; n16715
g16460 and n16714_not n16715_not ; n16716
g16461 and n16615_not n16716 ; n16717
g16462 and n16716 n16717_not ; n16718
g16463 and n16615_not n16717_not ; n16719
g16464 and n16718_not n16719_not ; n16720
g16465 and n16407_not n16420_not ; n16721
g16466 and n16720 n16721 ; n16722
g16467 and n16720_not n16721_not ; n16723
g16468 and n16722_not n16723_not ; n16724
g16469 and b[29] n6595 ; n16725
g16470 and b[27] n6902 ; n16726
g16471 and b[28] n6590 ; n16727
g16472 and n16726_not n16727_not ; n16728
g16473 and n16725_not n16728 ; n16729
g16474 and n3383 n6598 ; n16730
g16475 and n16729 n16730_not ; n16731
g16476 and a[44] n16731_not ; n16732
g16477 and a[44] n16732_not ; n16733
g16478 and n16731_not n16732_not ; n16734
g16479 and n16733_not n16734_not ; n16735
g16480 and n16724 n16735_not ; n16736
g16481 and n16724 n16736_not ; n16737
g16482 and n16735_not n16736_not ; n16738
g16483 and n16737_not n16738_not ; n16739
g16484 and n16426_not n16439_not ; n16740
g16485 and n16739 n16740 ; n16741
g16486 and n16739_not n16740_not ; n16742
g16487 and n16741_not n16742_not ; n16743
g16488 and b[32] n5777 ; n16744
g16489 and b[30] n6059 ; n16745
g16490 and b[31] n5772 ; n16746
g16491 and n16745_not n16746_not ; n16747
g16492 and n16744_not n16747 ; n16748
g16493 and n4013 n5780 ; n16749
g16494 and n16748 n16749_not ; n16750
g16495 and a[41] n16750_not ; n16751
g16496 and a[41] n16751_not ; n16752
g16497 and n16750_not n16751_not ; n16753
g16498 and n16752_not n16753_not ; n16754
g16499 and n16743_not n16754 ; n16755
g16500 and n16743 n16754_not ; n16756
g16501 and n16755_not n16756_not ; n16757
g16502 and n16445_not n16459_not ; n16758
g16503 and n16757 n16758_not ; n16759
g16504 and n16757_not n16758 ; n16760
g16505 and n16759_not n16760_not ; n16761
g16506 and n16604_not n16761 ; n16762
g16507 and n16761 n16762_not ; n16763
g16508 and n16604_not n16762_not ; n16764
g16509 and n16763_not n16764_not ; n16765
g16510 and n16461_not n16464_not ; n16766
g16511 and n16765 n16766 ; n16767
g16512 and n16765_not n16766_not ; n16768
g16513 and n16767_not n16768_not ; n16769
g16514 and b[38] n4287 ; n16770
g16515 and b[36] n4532 ; n16771
g16516 and b[37] n4282 ; n16772
g16517 and n16771_not n16772_not ; n16773
g16518 and n16770_not n16773 ; n16774
g16519 and n4290 n5205 ; n16775
g16520 and n16774 n16775_not ; n16776
g16521 and a[35] n16776_not ; n16777
g16522 and a[35] n16777_not ; n16778
g16523 and n16776_not n16777_not ; n16779
g16524 and n16778_not n16779_not ; n16780
g16525 and n16769 n16780_not ; n16781
g16526 and n16769_not n16780 ; n16782
g16527 and n16593 n16782_not ; n16783
g16528 and n16781_not n16783 ; n16784
g16529 and n16593 n16784_not ; n16785
g16530 and n16782_not n16784_not ; n16786
g16531 and n16781_not n16786 ; n16787
g16532 and n16785_not n16787_not ; n16788
g16533 and n16280_not n16474_not ; n16789
g16534 and b[44] n3050 ; n16790
g16535 and b[42] n3243 ; n16791
g16536 and b[43] n3045 ; n16792
g16537 and n16791_not n16792_not ; n16793
g16538 and n16790_not n16793 ; n16794
g16539 and n3053_not n16794 ; n16795
g16540 and n7072_not n16794 ; n16796
g16541 and n16795_not n16796_not ; n16797
g16542 and a[29] n16797_not ; n16798
g16543 and a[29]_not n16797 ; n16799
g16544 and n16798_not n16799_not ; n16800
g16545 and n16789_not n16800_not ; n16801
g16546 and n16789_not n16801_not ; n16802
g16547 and n16800_not n16801_not ; n16803
g16548 and n16802_not n16803_not ; n16804
g16549 and n16788_not n16804_not ; n16805
g16550 and n16788_not n16805_not ; n16806
g16551 and n16804_not n16805_not ; n16807
g16552 and n16806_not n16807_not ; n16808
g16553 and n16578_not n16808_not ; n16809
g16554 and n16578_not n16809_not ; n16810
g16555 and n16808_not n16809_not ; n16811
g16556 and n16810_not n16811_not ; n16812
g16557 and n16561_not n16812 ; n16813
g16558 and n16561 n16812_not ; n16814
g16559 and n16813_not n16814_not ; n16815
g16560 and n16235_not n16484_not ; n16816
g16561 and n16232_not n16816_not ; n16817
g16562 and b[53] n1627 ; n16818
g16563 and b[51] n1763 ; n16819
g16564 and b[52] n1622 ; n16820
g16565 and n16819_not n16820_not ; n16821
g16566 and n16818_not n16821 ; n16822
g16567 and n1630_not n16822 ; n16823
g16568 and n9972_not n16822 ; n16824
g16569 and n16823_not n16824_not ; n16825
g16570 and a[20] n16825_not ; n16826
g16571 and a[20]_not n16825 ; n16827
g16572 and n16826_not n16827_not ; n16828
g16573 and n16817_not n16828_not ; n16829
g16574 and n16817_not n16829_not ; n16830
g16575 and n16828_not n16829_not ; n16831
g16576 and n16830_not n16831_not ; n16832
g16577 and n16815 n16832_not ; n16833
g16578 and n16815 n16833_not ; n16834
g16579 and n16832_not n16833_not ; n16835
g16580 and n16834_not n16835_not ; n16836
g16581 and n16546 n16836_not ; n16837
g16582 and n16546 n16837_not ; n16838
g16583 and n16836_not n16837_not ; n16839
g16584 and n16838_not n16839_not ; n16840
g16585 and b[59] n951 ; n16841
g16586 and b[57] n1056 ; n16842
g16587 and b[58] n946 ; n16843
g16588 and n16842_not n16843_not ; n16844
g16589 and n16841_not n16844 ; n16845
g16590 and n954 n12179 ; n16846
g16591 and n16845 n16846_not ; n16847
g16592 and a[14] n16847_not ; n16848
g16593 and a[14] n16848_not ; n16849
g16594 and n16847_not n16848_not ; n16850
g16595 and n16849_not n16850_not ; n16851
g16596 and n16202_not n16492_not ; n16852
g16597 and n16851_not n16852_not ; n16853
g16598 and n16851_not n16853_not ; n16854
g16599 and n16852_not n16853_not ; n16855
g16600 and n16854_not n16855_not ; n16856
g16601 and n16840_not n16856 ; n16857
g16602 and n16840 n16856_not ; n16858
g16603 and n16857_not n16858_not ; n16859
g16604 and n16186_not n16495_not ; n16860
g16605 and b[62] n700 ; n16861
g16606 and b[60] n767 ; n16862
g16607 and b[61] n695 ; n16863
g16608 and n16862_not n16863_not ; n16864
g16609 and n16861_not n16864 ; n16865
g16610 and n703_not n16865 ; n16866
g16611 and n13370_not n16865 ; n16867
g16612 and n16866_not n16867_not ; n16868
g16613 and a[11] n16868_not ; n16869
g16614 and a[11]_not n16868 ; n16870
g16615 and n16869_not n16870_not ; n16871
g16616 and n16860_not n16871_not ; n16872
g16617 and n16860_not n16872_not ; n16873
g16618 and n16871_not n16872_not ; n16874
g16619 and n16873_not n16874_not ; n16875
g16620 and n16859_not n16875_not ; n16876
g16621 and n16859 n16874_not ; n16877
g16622 and n16873_not n16877 ; n16878
g16623 and n16876_not n16878_not ; n16879
g16624 and n16531_not n16879 ; n16880
g16625 and n16531 n16879_not ; n16881
g16626 and n16880_not n16881_not ; n16882
g16627 and n16519_not n16882 ; n16883
g16628 and n16519_not n16883_not ; n16884
g16629 and n16882 n16883_not ; n16885
g16630 and n16884_not n16885_not ; n16886
g16631 and n16518_not n16886_not ; n16887
g16632 and n16518 n16885_not ; n16888
g16633 and n16884_not n16888 ; n16889
g16634 and n16887_not n16889_not ; f[71]
g16635 and n16883_not n16887_not ; n16891
g16636 and n16528_not n16880_not ; n16892
g16637 and n16872_not n16876_not ; n16893
g16638 and b[63] n700 ; n16894
g16639 and b[61] n767 ; n16895
g16640 and b[62] n695 ; n16896
g16641 and n16895_not n16896_not ; n16897
g16642 and n16894_not n16897 ; n16898
g16643 and n703 n13771 ; n16899
g16644 and n16898 n16899_not ; n16900
g16645 and a[11] n16900_not ; n16901
g16646 and a[11] n16901_not ; n16902
g16647 and n16900_not n16901_not ; n16903
g16648 and n16902_not n16903_not ; n16904
g16649 and n16893_not n16904_not ; n16905
g16650 and n16893_not n16905_not ; n16906
g16651 and n16904_not n16905_not ; n16907
g16652 and n16906_not n16907_not ; n16908
g16653 and n16840_not n16856_not ; n16909
g16654 and n16853_not n16909_not ; n16910
g16655 and b[60] n951 ; n16911
g16656 and b[58] n1056 ; n16912
g16657 and b[59] n946 ; n16913
g16658 and n16912_not n16913_not ; n16914
g16659 and n16911_not n16914 ; n16915
g16660 and n954 n12211 ; n16916
g16661 and n16915 n16916_not ; n16917
g16662 and a[14] n16917_not ; n16918
g16663 and a[14] n16918_not ; n16919
g16664 and n16917_not n16918_not ; n16920
g16665 and n16919_not n16920_not ; n16921
g16666 and n16910_not n16921 ; n16922
g16667 and n16910 n16921_not ; n16923
g16668 and n16922_not n16923_not ; n16924
g16669 and b[57] n1302 ; n16925
g16670 and b[55] n1391 ; n16926
g16671 and b[56] n1297 ; n16927
g16672 and n16926_not n16927_not ; n16928
g16673 and n16925_not n16928 ; n16929
g16674 and n1305 n11410 ; n16930
g16675 and n16929 n16930_not ; n16931
g16676 and a[17] n16931_not ; n16932
g16677 and a[17] n16932_not ; n16933
g16678 and n16931_not n16932_not ; n16934
g16679 and n16933_not n16934_not ; n16935
g16680 and n16545_not n16837_not ; n16936
g16681 and n16935 n16936 ; n16937
g16682 and n16935_not n16936_not ; n16938
g16683 and n16937_not n16938_not ; n16939
g16684 and n16829_not n16833_not ; n16940
g16685 and b[54] n1627 ; n16941
g16686 and b[52] n1763 ; n16942
g16687 and b[53] n1622 ; n16943
g16688 and n16942_not n16943_not ; n16944
g16689 and n16941_not n16944 ; n16945
g16690 and n1630 n9998 ; n16946
g16691 and n16945 n16946_not ; n16947
g16692 and a[20] n16947_not ; n16948
g16693 and a[20] n16948_not ; n16949
g16694 and n16947_not n16948_not ; n16950
g16695 and n16949_not n16950_not ; n16951
g16696 and n16940_not n16951_not ; n16952
g16697 and n16940_not n16952_not ; n16953
g16698 and n16951_not n16952_not ; n16954
g16699 and n16953_not n16954_not ; n16955
g16700 and b[48] n2539 ; n16956
g16701 and b[46] n2685 ; n16957
g16702 and b[47] n2534 ; n16958
g16703 and n16957_not n16958_not ; n16959
g16704 and n16956_not n16959 ; n16960
g16705 and n2542 n8009 ; n16961
g16706 and n16960 n16961_not ; n16962
g16707 and a[26] n16962_not ; n16963
g16708 and a[26] n16963_not ; n16964
g16709 and n16962_not n16963_not ; n16965
g16710 and n16964_not n16965_not ; n16966
g16711 and n16575_not n16809_not ; n16967
g16712 and n16966 n16967 ; n16968
g16713 and n16966_not n16967_not ; n16969
g16714 and n16968_not n16969_not ; n16970
g16715 and n16801_not n16805_not ; n16971
g16716 and b[45] n3050 ; n16972
g16717 and b[43] n3243 ; n16973
g16718 and b[44] n3045 ; n16974
g16719 and n16973_not n16974_not ; n16975
g16720 and n16972_not n16975 ; n16976
g16721 and n3053 n7361 ; n16977
g16722 and n16976 n16977_not ; n16978
g16723 and a[29] n16978_not ; n16979
g16724 and a[29] n16979_not ; n16980
g16725 and n16978_not n16979_not ; n16981
g16726 and n16980_not n16981_not ; n16982
g16727 and n16971_not n16982_not ; n16983
g16728 and n16971_not n16983_not ; n16984
g16729 and n16982_not n16983_not ; n16985
g16730 and n16984_not n16985_not ; n16986
g16731 and n16592_not n16784_not ; n16987
g16732 and b[42] n3638 ; n16988
g16733 and b[40] n3843 ; n16989
g16734 and b[41] n3633 ; n16990
g16735 and n16989_not n16990_not ; n16991
g16736 and n16988_not n16991 ; n16992
g16737 and n3641 n6489 ; n16993
g16738 and n16992 n16993_not ; n16994
g16739 and a[32] n16994_not ; n16995
g16740 and a[32] n16995_not ; n16996
g16741 and n16994_not n16995_not ; n16997
g16742 and n16996_not n16997_not ; n16998
g16743 and n16987_not n16998_not ; n16999
g16744 and n16987_not n16999_not ; n17000
g16745 and n16998_not n16999_not ; n17001
g16746 and n17000_not n17001_not ; n17002
g16747 and n16759_not n16762_not ; n17003
g16748 and n16742_not n16756_not ; n17004
g16749 and n16723_not n16736_not ; n17005
g16750 and n16706_not n16710_not ; n17006
g16751 and b[24] n8362 ; n17007
g16752 and b[22] n8715 ; n17008
g16753 and b[23] n8357 ; n17009
g16754 and n17008_not n17009_not ; n17010
g16755 and n17007_not n17010 ; n17011
g16756 and n2458 n8365 ; n17012
g16757 and n17011 n17012_not ; n17013
g16758 and a[50] n17013_not ; n17014
g16759 and a[50] n17014_not ; n17015
g16760 and n17013_not n17014_not ; n17016
g16761 and n17015_not n17016_not ; n17017
g16762 and b[18] n10426 ; n17018
g16763 and b[16] n10796 ; n17019
g16764 and b[17] n10421 ; n17020
g16765 and n17019_not n17020_not ; n17021
g16766 and n17018_not n17021 ; n17022
g16767 and n1566 n10429 ; n17023
g16768 and n17022 n17023_not ; n17024
g16769 and a[56] n17024_not ; n17025
g16770 and a[56] n17025_not ; n17026
g16771 and n17024_not n17025_not ; n17027
g16772 and n17026_not n17027_not ; n17028
g16773 and n16641_not n16652_not ; n17029
g16774 and n16667_not n17029_not ; n17030
g16775 and b[12] n12668 ; n17031
g16776 and b[10] n13047 ; n17032
g16777 and b[11] n12663 ; n17033
g16778 and n17032_not n17033_not ; n17034
g16779 and n17031_not n17034 ; n17035
g16780 and n842 n12671 ; n17036
g16781 and n17035 n17036_not ; n17037
g16782 and a[62] n17037_not ; n17038
g16783 and a[62] n17038_not ; n17039
g16784 and n17037_not n17038_not ; n17040
g16785 and n17039_not n17040_not ; n17041
g16786 and b[8] n13903 ; n17042
g16787 and b[9] n13488_not ; n17043
g16788 and n17042_not n17043_not ; n17044
g16789 and a[8] n16633_not ; n17045
g16790 and a[8]_not n16633 ; n17046
g16791 and n17045_not n17046_not ; n17047
g16792 and n17044_not n17047_not ; n17048
g16793 and n17044 n17047 ; n17049
g16794 and n17048_not n17049_not ; n17050
g16795 and n16639_not n17050 ; n17051
g16796 and n16639 n17050_not ; n17052
g16797 and n17051_not n17052_not ; n17053
g16798 and n17041 n17053 ; n17054
g16799 and n17041_not n17053_not ; n17055
g16800 and n17054_not n17055_not ; n17056
g16801 and b[15] n11531 ; n17057
g16802 and b[13] n11896 ; n17058
g16803 and b[14] n11526 ; n17059
g16804 and n17058_not n17059_not ; n17060
g16805 and n17057_not n17060 ; n17061
g16806 and n1131 n11534 ; n17062
g16807 and n17061 n17062_not ; n17063
g16808 and a[59] n17063_not ; n17064
g16809 and a[59] n17064_not ; n17065
g16810 and n17063_not n17064_not ; n17066
g16811 and n17065_not n17066_not ; n17067
g16812 and n17056_not n17067_not ; n17068
g16813 and n17056 n17067 ; n17069
g16814 and n17068_not n17069_not ; n17070
g16815 and n17030_not n17070 ; n17071
g16816 and n17030 n17070_not ; n17072
g16817 and n17071_not n17072_not ; n17073
g16818 and n17028_not n17073 ; n17074
g16819 and n17073 n17074_not ; n17075
g16820 and n17028_not n17074_not ; n17076
g16821 and n17075_not n17076_not ; n17077
g16822 and n16671_not n16684_not ; n17078
g16823 and n17077 n17078 ; n17079
g16824 and n17077_not n17078_not ; n17080
g16825 and n17079_not n17080_not ; n17081
g16826 and b[21] n9339 ; n17082
g16827 and b[19] n9732 ; n17083
g16828 and b[20] n9334 ; n17084
g16829 and n17083_not n17084_not ; n17085
g16830 and n17082_not n17085 ; n17086
g16831 and n1984 n9342 ; n17087
g16832 and n17086 n17087_not ; n17088
g16833 and a[53] n17088_not ; n17089
g16834 and a[53] n17089_not ; n17090
g16835 and n17088_not n17089_not ; n17091
g16836 and n17090_not n17091_not ; n17092
g16837 and n17081 n17092_not ; n17093
g16838 and n17081 n17093_not ; n17094
g16839 and n17092_not n17093_not ; n17095
g16840 and n17094_not n17095_not ; n17096
g16841 and n16690_not n16704_not ; n17097
g16842 and n17096_not n17097_not ; n17098
g16843 and n17096 n17097 ; n17099
g16844 and n17098_not n17099_not ; n17100
g16845 and n17017_not n17100 ; n17101
g16846 and n17017_not n17101_not ; n17102
g16847 and n17100 n17101_not ; n17103
g16848 and n17102_not n17103_not ; n17104
g16849 and n17006_not n17104_not ; n17105
g16850 and n17006_not n17105_not ; n17106
g16851 and n17104_not n17105_not ; n17107
g16852 and n17106_not n17107_not ; n17108
g16853 and b[27] n7446 ; n17109
g16854 and b[25] n7787 ; n17110
g16855 and b[26] n7441 ; n17111
g16856 and n17110_not n17111_not ; n17112
g16857 and n17109_not n17112 ; n17113
g16858 and n2990 n7449 ; n17114
g16859 and n17113 n17114_not ; n17115
g16860 and a[47] n17115_not ; n17116
g16861 and a[47] n17116_not ; n17117
g16862 and n17115_not n17116_not ; n17118
g16863 and n17117_not n17118_not ; n17119
g16864 and n17108_not n17119_not ; n17120
g16865 and n17108_not n17120_not ; n17121
g16866 and n17119_not n17120_not ; n17122
g16867 and n17121_not n17122_not ; n17123
g16868 and n16714_not n16717_not ; n17124
g16869 and n17123 n17124 ; n17125
g16870 and n17123_not n17124_not ; n17126
g16871 and n17125_not n17126_not ; n17127
g16872 and b[30] n6595 ; n17128
g16873 and b[28] n6902 ; n17129
g16874 and b[29] n6590 ; n17130
g16875 and n17129_not n17130_not ; n17131
g16876 and n17128_not n17131 ; n17132
g16877 and n3577 n6598 ; n17133
g16878 and n17132 n17133_not ; n17134
g16879 and a[44] n17134_not ; n17135
g16880 and a[44] n17135_not ; n17136
g16881 and n17134_not n17135_not ; n17137
g16882 and n17136_not n17137_not ; n17138
g16883 and n17127 n17138_not ; n17139
g16884 and n17127_not n17138 ; n17140
g16885 and n17005_not n17140_not ; n17141
g16886 and n17139_not n17141 ; n17142
g16887 and n17005_not n17142_not ; n17143
g16888 and n17139_not n17142_not ; n17144
g16889 and n17140_not n17144 ; n17145
g16890 and n17143_not n17145_not ; n17146
g16891 and b[33] n5777 ; n17147
g16892 and b[31] n6059 ; n17148
g16893 and b[32] n5772 ; n17149
g16894 and n17148_not n17149_not ; n17150
g16895 and n17147_not n17150 ; n17151
g16896 and n4223 n5780 ; n17152
g16897 and n17151 n17152_not ; n17153
g16898 and a[41] n17153_not ; n17154
g16899 and a[41] n17154_not ; n17155
g16900 and n17153_not n17154_not ; n17156
g16901 and n17155_not n17156_not ; n17157
g16902 and n17146_not n17157_not ; n17158
g16903 and n17146_not n17158_not ; n17159
g16904 and n17157_not n17158_not ; n17160
g16905 and n17159_not n17160_not ; n17161
g16906 and n17004_not n17161 ; n17162
g16907 and n17004 n17161_not ; n17163
g16908 and n17162_not n17163_not ; n17164
g16909 and b[36] n5035 ; n17165
g16910 and b[34] n5277 ; n17166
g16911 and b[35] n5030 ; n17167
g16912 and n17166_not n17167_not ; n17168
g16913 and n17165_not n17168 ; n17169
g16914 and n4922 n5038 ; n17170
g16915 and n17169 n17170_not ; n17171
g16916 and a[38] n17171_not ; n17172
g16917 and a[38] n17172_not ; n17173
g16918 and n17171_not n17172_not ; n17174
g16919 and n17173_not n17174_not ; n17175
g16920 and n17164_not n17175_not ; n17176
g16921 and n17164 n17175 ; n17177
g16922 and n17176_not n17177_not ; n17178
g16923 and n17003 n17178_not ; n17179
g16924 and n17003_not n17178 ; n17180
g16925 and n17179_not n17180_not ; n17181
g16926 and b[39] n4287 ; n17182
g16927 and b[37] n4532 ; n17183
g16928 and b[38] n4282 ; n17184
g16929 and n17183_not n17184_not ; n17185
g16930 and n17182_not n17185 ; n17186
g16931 and n4290 n5451 ; n17187
g16932 and n17186 n17187_not ; n17188
g16933 and a[35] n17188_not ; n17189
g16934 and a[35] n17189_not ; n17190
g16935 and n17188_not n17189_not ; n17191
g16936 and n17190_not n17191_not ; n17192
g16937 and n17181 n17192_not ; n17193
g16938 and n17181 n17193_not ; n17194
g16939 and n17192_not n17193_not ; n17195
g16940 and n17194_not n17195_not ; n17196
g16941 and n16768_not n16781_not ; n17197
g16942 and n17196_not n17197_not ; n17198
g16943 and n17196_not n17198_not ; n17199
g16944 and n17197_not n17198_not ; n17200
g16945 and n17199_not n17200_not ; n17201
g16946 and n17002_not n17201_not ; n17202
g16947 and n17002_not n17202_not ; n17203
g16948 and n17201_not n17202_not ; n17204
g16949 and n17203_not n17204_not ; n17205
g16950 and n16986_not n17205 ; n17206
g16951 and n16986 n17205_not ; n17207
g16952 and n17206_not n17207_not ; n17208
g16953 and n16970 n17208_not ; n17209
g16954 and n16970 n17209_not ; n17210
g16955 and n17208_not n17209_not ; n17211
g16956 and n17210_not n17211_not ; n17212
g16957 and b[51] n2048 ; n17213
g16958 and b[49] n2198 ; n17214
g16959 and b[50] n2043 ; n17215
g16960 and n17214_not n17215_not ; n17216
g16961 and n17213_not n17216 ; n17217
g16962 and n2051 n8976 ; n17218
g16963 and n17217 n17218_not ; n17219
g16964 and a[23] n17219_not ; n17220
g16965 and a[23] n17220_not ; n17221
g16966 and n17219_not n17220_not ; n17222
g16967 and n17221_not n17222_not ; n17223
g16968 and n16560_not n16814_not ; n17224
g16969 and n17223_not n17224_not ; n17225
g16970 and n17223 n17224 ; n17226
g16971 and n17225_not n17226_not ; n17227
g16972 and n17212_not n17227 ; n17228
g16973 and n17212_not n17228_not ; n17229
g16974 and n17227 n17228_not ; n17230
g16975 and n17229_not n17230_not ; n17231
g16976 and n16955_not n17231_not ; n17232
g16977 and n16955_not n17232_not ; n17233
g16978 and n17231_not n17232_not ; n17234
g16979 and n17233_not n17234_not ; n17235
g16980 and n16939 n17235_not ; n17236
g16981 and n16939_not n17235 ; n17237
g16982 and n16924_not n17237_not ; n17238
g16983 and n17236_not n17238 ; n17239
g16984 and n16924_not n17239_not ; n17240
g16985 and n17237_not n17239_not ; n17241
g16986 and n17236_not n17241 ; n17242
g16987 and n17240_not n17242_not ; n17243
g16988 and n16908_not n17243 ; n17244
g16989 and n16908 n17243_not ; n17245
g16990 and n17244_not n17245_not ; n17246
g16991 and n16892_not n17246_not ; n17247
g16992 and n16892_not n17247_not ; n17248
g16993 and n17246_not n17247_not ; n17249
g16994 and n17248_not n17249_not ; n17250
g16995 and n16891_not n17250_not ; n17251
g16996 and n16891 n17249_not ; n17252
g16997 and n17248_not n17252 ; n17253
g16998 and n17251_not n17253_not ; f[72]
g16999 and n17247_not n17251_not ; n17255
g17000 and n16908_not n17243_not ; n17256
g17001 and n16905_not n17256_not ; n17257
g17002 and b[61] n951 ; n17258
g17003 and b[59] n1056 ; n17259
g17004 and b[60] n946 ; n17260
g17005 and n17259_not n17260_not ; n17261
g17006 and n17258_not n17261 ; n17262
g17007 and n954 n12969 ; n17263
g17008 and n17262 n17263_not ; n17264
g17009 and a[14] n17264_not ; n17265
g17010 and a[14] n17265_not ; n17266
g17011 and n17264_not n17265_not ; n17267
g17012 and n17266_not n17267_not ; n17268
g17013 and n16938_not n17236_not ; n17269
g17014 and n17268_not n17269_not ; n17270
g17015 and n17268_not n17270_not ; n17271
g17016 and n17269_not n17270_not ; n17272
g17017 and n17271_not n17272_not ; n17273
g17018 and b[55] n1627 ; n17274
g17019 and b[53] n1763 ; n17275
g17020 and b[54] n1622 ; n17276
g17021 and n17275_not n17276_not ; n17277
g17022 and n17274_not n17277 ; n17278
g17023 and n1630 n10684 ; n17279
g17024 and n17278 n17279_not ; n17280
g17025 and a[20] n17280_not ; n17281
g17026 and a[20] n17281_not ; n17282
g17027 and n17280_not n17281_not ; n17283
g17028 and n17282_not n17283_not ; n17284
g17029 and n17225_not n17228_not ; n17285
g17030 and n17284 n17285 ; n17286
g17031 and n17284_not n17285_not ; n17287
g17032 and n17286_not n17287_not ; n17288
g17033 and b[52] n2048 ; n17289
g17034 and b[50] n2198 ; n17290
g17035 and b[51] n2043 ; n17291
g17036 and n17290_not n17291_not ; n17292
g17037 and n17289_not n17292 ; n17293
g17038 and n2051 n9628 ; n17294
g17039 and n17293 n17294_not ; n17295
g17040 and a[23] n17295_not ; n17296
g17041 and a[23] n17296_not ; n17297
g17042 and n17295_not n17296_not ; n17298
g17043 and n17297_not n17298_not ; n17299
g17044 and n16969_not n17209_not ; n17300
g17045 and n17299 n17300 ; n17301
g17046 and n17299_not n17300_not ; n17302
g17047 and n17301_not n17302_not ; n17303
g17048 and b[49] n2539 ; n17304
g17049 and b[47] n2685 ; n17305
g17050 and b[48] n2534 ; n17306
g17051 and n17305_not n17306_not ; n17307
g17052 and n17304_not n17307 ; n17308
g17053 and n2542 n8625 ; n17309
g17054 and n17308 n17309_not ; n17310
g17055 and a[26] n17310_not ; n17311
g17056 and a[26] n17311_not ; n17312
g17057 and n17310_not n17311_not ; n17313
g17058 and n17312_not n17313_not ; n17314
g17059 and n16986_not n17205_not ; n17315
g17060 and n16983_not n17315_not ; n17316
g17061 and n17314_not n17316_not ; n17317
g17062 and n17314_not n17317_not ; n17318
g17063 and n17316_not n17317_not ; n17319
g17064 and n17318_not n17319_not ; n17320
g17065 and b[43] n3638 ; n17321
g17066 and b[41] n3843 ; n17322
g17067 and b[42] n3633 ; n17323
g17068 and n17322_not n17323_not ; n17324
g17069 and n17321_not n17324 ; n17325
g17070 and n3641 n6515 ; n17326
g17071 and n17325 n17326_not ; n17327
g17072 and a[32] n17327_not ; n17328
g17073 and a[32] n17328_not ; n17329
g17074 and n17327_not n17328_not ; n17330
g17075 and n17329_not n17330_not ; n17331
g17076 and n17193_not n17198_not ; n17332
g17077 and n17331 n17332 ; n17333
g17078 and n17331_not n17332_not ; n17334
g17079 and n17333_not n17334_not ; n17335
g17080 and b[40] n4287 ; n17336
g17081 and b[38] n4532 ; n17337
g17082 and b[39] n4282 ; n17338
g17083 and n17337_not n17338_not ; n17339
g17084 and n17336_not n17339 ; n17340
g17085 and n4290 n5955 ; n17341
g17086 and n17340 n17341_not ; n17342
g17087 and a[35] n17342_not ; n17343
g17088 and a[35] n17343_not ; n17344
g17089 and n17342_not n17343_not ; n17345
g17090 and n17344_not n17345_not ; n17346
g17091 and n17176_not n17180_not ; n17347
g17092 and b[37] n5035 ; n17348
g17093 and b[35] n5277 ; n17349
g17094 and b[36] n5030 ; n17350
g17095 and n17349_not n17350_not ; n17351
g17096 and n17348_not n17351 ; n17352
g17097 and n5038 n5181 ; n17353
g17098 and n17352 n17353_not ; n17354
g17099 and a[38] n17354_not ; n17355
g17100 and a[38] n17355_not ; n17356
g17101 and n17354_not n17355_not ; n17357
g17102 and n17356_not n17357_not ; n17358
g17103 and n17004_not n17161_not ; n17359
g17104 and n17158_not n17359_not ; n17360
g17105 and b[34] n5777 ; n17361
g17106 and b[32] n6059 ; n17362
g17107 and b[33] n5772 ; n17363
g17108 and n17362_not n17363_not ; n17364
g17109 and n17361_not n17364 ; n17365
g17110 and n4466 n5780 ; n17366
g17111 and n17365 n17366_not ; n17367
g17112 and a[41] n17367_not ; n17368
g17113 and a[41] n17368_not ; n17369
g17114 and n17367_not n17368_not ; n17370
g17115 and n17369_not n17370_not ; n17371
g17116 and b[13] n12668 ; n17372
g17117 and b[11] n13047 ; n17373
g17118 and b[12] n12663 ; n17374
g17119 and n17373_not n17374_not ; n17375
g17120 and n17372_not n17375 ; n17376
g17121 and n1008 n12671 ; n17377
g17122 and n17376 n17377_not ; n17378
g17123 and a[62] n17378_not ; n17379
g17124 and a[62] n17379_not ; n17380
g17125 and n17378_not n17379_not ; n17381
g17126 and n17380_not n17381_not ; n17382
g17127 and b[9] n13903 ; n17383
g17128 and b[10] n13488_not ; n17384
g17129 and n17383_not n17384_not ; n17385
g17130 and a[8]_not n16633_not ; n17386
g17131 and n17048_not n17386_not ; n17387
g17132 and n17385 n17387_not ; n17388
g17133 and n17385 n17388_not ; n17389
g17134 and n17387_not n17388_not ; n17390
g17135 and n17389_not n17390_not ; n17391
g17136 and n17382_not n17391_not ; n17392
g17137 and n17382_not n17392_not ; n17393
g17138 and n17391_not n17392_not ; n17394
g17139 and n17393_not n17394_not ; n17395
g17140 and n17041_not n17053 ; n17396
g17141 and n17051_not n17396_not ; n17397
g17142 and n17395_not n17397_not ; n17398
g17143 and n17395_not n17398_not ; n17399
g17144 and n17397_not n17398_not ; n17400
g17145 and n17399_not n17400_not ; n17401
g17146 and b[16] n11531 ; n17402
g17147 and b[14] n11896 ; n17403
g17148 and b[15] n11526 ; n17404
g17149 and n17403_not n17404_not ; n17405
g17150 and n17402_not n17405 ; n17406
g17151 and n1237 n11534 ; n17407
g17152 and n17406 n17407_not ; n17408
g17153 and a[59] n17408_not ; n17409
g17154 and a[59] n17409_not ; n17410
g17155 and n17408_not n17409_not ; n17411
g17156 and n17410_not n17411_not ; n17412
g17157 and n17401_not n17412_not ; n17413
g17158 and n17401_not n17413_not ; n17414
g17159 and n17412_not n17413_not ; n17415
g17160 and n17414_not n17415_not ; n17416
g17161 and n17068_not n17071_not ; n17417
g17162 and n17416 n17417 ; n17418
g17163 and n17416_not n17417_not ; n17419
g17164 and n17418_not n17419_not ; n17420
g17165 and b[19] n10426 ; n17421
g17166 and b[17] n10796 ; n17422
g17167 and b[18] n10421 ; n17423
g17168 and n17422_not n17423_not ; n17424
g17169 and n17421_not n17424 ; n17425
g17170 and n1708 n10429 ; n17426
g17171 and n17425 n17426_not ; n17427
g17172 and a[56] n17427_not ; n17428
g17173 and a[56] n17428_not ; n17429
g17174 and n17427_not n17428_not ; n17430
g17175 and n17429_not n17430_not ; n17431
g17176 and n17420 n17431_not ; n17432
g17177 and n17420 n17432_not ; n17433
g17178 and n17431_not n17432_not ; n17434
g17179 and n17433_not n17434_not ; n17435
g17180 and n17074_not n17080_not ; n17436
g17181 and n17435 n17436 ; n17437
g17182 and n17435_not n17436_not ; n17438
g17183 and n17437_not n17438_not ; n17439
g17184 and b[22] n9339 ; n17440
g17185 and b[20] n9732 ; n17441
g17186 and b[21] n9334 ; n17442
g17187 and n17441_not n17442_not ; n17443
g17188 and n17440_not n17443 ; n17444
g17189 and n2145 n9342 ; n17445
g17190 and n17444 n17445_not ; n17446
g17191 and a[53] n17446_not ; n17447
g17192 and a[53] n17447_not ; n17448
g17193 and n17446_not n17447_not ; n17449
g17194 and n17448_not n17449_not ; n17450
g17195 and n17439 n17450_not ; n17451
g17196 and n17439 n17451_not ; n17452
g17197 and n17450_not n17451_not ; n17453
g17198 and n17452_not n17453_not ; n17454
g17199 and n17093_not n17098_not ; n17455
g17200 and n17454 n17455 ; n17456
g17201 and n17454_not n17455_not ; n17457
g17202 and n17456_not n17457_not ; n17458
g17203 and b[25] n8362 ; n17459
g17204 and b[23] n8715 ; n17460
g17205 and b[24] n8357 ; n17461
g17206 and n17460_not n17461_not ; n17462
g17207 and n17459_not n17462 ; n17463
g17208 and n2485 n8365 ; n17464
g17209 and n17463 n17464_not ; n17465
g17210 and a[50] n17465_not ; n17466
g17211 and a[50] n17466_not ; n17467
g17212 and n17465_not n17466_not ; n17468
g17213 and n17467_not n17468_not ; n17469
g17214 and n17458 n17469_not ; n17470
g17215 and n17458 n17470_not ; n17471
g17216 and n17469_not n17470_not ; n17472
g17217 and n17471_not n17472_not ; n17473
g17218 and n17101_not n17105_not ; n17474
g17219 and n17473 n17474 ; n17475
g17220 and n17473_not n17474_not ; n17476
g17221 and n17475_not n17476_not ; n17477
g17222 and b[28] n7446 ; n17478
g17223 and b[26] n7787 ; n17479
g17224 and b[27] n7441 ; n17480
g17225 and n17479_not n17480_not ; n17481
g17226 and n17478_not n17481 ; n17482
g17227 and n3189 n7449 ; n17483
g17228 and n17482 n17483_not ; n17484
g17229 and a[47] n17484_not ; n17485
g17230 and a[47] n17485_not ; n17486
g17231 and n17484_not n17485_not ; n17487
g17232 and n17486_not n17487_not ; n17488
g17233 and n17477 n17488_not ; n17489
g17234 and n17477 n17489_not ; n17490
g17235 and n17488_not n17489_not ; n17491
g17236 and n17490_not n17491_not ; n17492
g17237 and n17120_not n17126_not ; n17493
g17238 and n17492 n17493 ; n17494
g17239 and n17492_not n17493_not ; n17495
g17240 and n17494_not n17495_not ; n17496
g17241 and b[31] n6595 ; n17497
g17242 and b[29] n6902 ; n17498
g17243 and b[30] n6590 ; n17499
g17244 and n17498_not n17499_not ; n17500
g17245 and n17497_not n17500 ; n17501
g17246 and n3796 n6598 ; n17502
g17247 and n17501 n17502_not ; n17503
g17248 and a[44] n17503_not ; n17504
g17249 and a[44] n17504_not ; n17505
g17250 and n17503_not n17504_not ; n17506
g17251 and n17505_not n17506_not ; n17507
g17252 and n17496_not n17507 ; n17508
g17253 and n17496 n17507_not ; n17509
g17254 and n17508_not n17509_not ; n17510
g17255 and n17144_not n17510 ; n17511
g17256 and n17144 n17510_not ; n17512
g17257 and n17511_not n17512_not ; n17513
g17258 and n17371_not n17513 ; n17514
g17259 and n17371 n17513_not ; n17515
g17260 and n17514_not n17515_not ; n17516
g17261 and n17360_not n17516 ; n17517
g17262 and n17360_not n17517_not ; n17518
g17263 and n17516 n17517_not ; n17519
g17264 and n17518_not n17519_not ; n17520
g17265 and n17358_not n17520_not ; n17521
g17266 and n17358 n17519_not ; n17522
g17267 and n17518_not n17522 ; n17523
g17268 and n17521_not n17523_not ; n17524
g17269 and n17347_not n17524 ; n17525
g17270 and n17347_not n17525_not ; n17526
g17271 and n17524 n17525_not ; n17527
g17272 and n17526_not n17527_not ; n17528
g17273 and n17346_not n17528_not ; n17529
g17274 and n17346_not n17529_not ; n17530
g17275 and n17528_not n17529_not ; n17531
g17276 and n17530_not n17531_not ; n17532
g17277 and n17335 n17532_not ; n17533
g17278 and n17335 n17533_not ; n17534
g17279 and n17532_not n17533_not ; n17535
g17280 and n17534_not n17535_not ; n17536
g17281 and n16999_not n17202_not ; n17537
g17282 and b[46] n3050 ; n17538
g17283 and b[44] n3243 ; n17539
g17284 and b[45] n3045 ; n17540
g17285 and n17539_not n17540_not ; n17541
g17286 and n17538_not n17541 ; n17542
g17287 and n3053_not n17542 ; n17543
g17288 and n7677_not n17542 ; n17544
g17289 and n17543_not n17544_not ; n17545
g17290 and a[29] n17545_not ; n17546
g17291 and a[29]_not n17545 ; n17547
g17292 and n17546_not n17547_not ; n17548
g17293 and n17537_not n17548_not ; n17549
g17294 and n17537_not n17549_not ; n17550
g17295 and n17548_not n17549_not ; n17551
g17296 and n17550_not n17551_not ; n17552
g17297 and n17536_not n17552_not ; n17553
g17298 and n17536_not n17553_not ; n17554
g17299 and n17552_not n17553_not ; n17555
g17300 and n17554_not n17555_not ; n17556
g17301 and n17320_not n17556_not ; n17557
g17302 and n17320_not n17557_not ; n17558
g17303 and n17556_not n17557_not ; n17559
g17304 and n17558_not n17559_not ; n17560
g17305 and n17303 n17560_not ; n17561
g17306 and n17303_not n17560 ; n17562
g17307 and n17288 n17562_not ; n17563
g17308 and n17561_not n17563 ; n17564
g17309 and n17288 n17564_not ; n17565
g17310 and n17562_not n17564_not ; n17566
g17311 and n17561_not n17566 ; n17567
g17312 and n17565_not n17567_not ; n17568
g17313 and n16952_not n17232_not ; n17569
g17314 and b[58] n1302 ; n17570
g17315 and b[56] n1391 ; n17571
g17316 and b[57] n1297 ; n17572
g17317 and n17571_not n17572_not ; n17573
g17318 and n17570_not n17573 ; n17574
g17319 and n1305_not n17574 ; n17575
g17320 and n11436_not n17574 ; n17576
g17321 and n17575_not n17576_not ; n17577
g17322 and a[17] n17577_not ; n17578
g17323 and a[17]_not n17577 ; n17579
g17324 and n17578_not n17579_not ; n17580
g17325 and n17569_not n17580_not ; n17581
g17326 and n17569_not n17581_not ; n17582
g17327 and n17580_not n17581_not ; n17583
g17328 and n17582_not n17583_not ; n17584
g17329 and n17568_not n17584_not ; n17585
g17330 and n17568_not n17585_not ; n17586
g17331 and n17584_not n17585_not ; n17587
g17332 and n17586_not n17587_not ; n17588
g17333 and n17273_not n17588_not ; n17589
g17334 and n17273_not n17589_not ; n17590
g17335 and n17588_not n17589_not ; n17591
g17336 and n17590_not n17591_not ; n17592
g17337 and n16910_not n16921_not ; n17593
g17338 and n17239_not n17593_not ; n17594
g17339 and b[62] n767 ; n17595
g17340 and b[63] n695 ; n17596
g17341 and n17595_not n17596_not ; n17597
g17342 and n703_not n17597 ; n17598
g17343 and n13800 n17597 ; n17599
g17344 and n17598_not n17599_not ; n17600
g17345 and a[11] n17600_not ; n17601
g17346 and a[11]_not n17600 ; n17602
g17347 and n17601_not n17602_not ; n17603
g17348 and n17594_not n17603_not ; n17604
g17349 and n17594_not n17604_not ; n17605
g17350 and n17603_not n17604_not ; n17606
g17351 and n17605_not n17606_not ; n17607
g17352 and n17592_not n17607_not ; n17608
g17353 and n17592 n17606_not ; n17609
g17354 and n17605_not n17609 ; n17610
g17355 and n17608_not n17610_not ; n17611
g17356 and n17257_not n17611 ; n17612
g17357 and n17257_not n17612_not ; n17613
g17358 and n17611 n17612_not ; n17614
g17359 and n17613_not n17614_not ; n17615
g17360 and n17255_not n17615_not ; n17616
g17361 and n17255 n17614_not ; n17617
g17362 and n17613_not n17617 ; n17618
g17363 and n17616_not n17618_not ; f[73]
g17364 and n17612_not n17616_not ; n17620
g17365 and n17604_not n17608_not ; n17621
g17366 and n17270_not n17589_not ; n17622
g17367 and b[63] n767 ; n17623
g17368 and n703 n13797 ; n17624
g17369 and n17623_not n17624_not ; n17625
g17370 and a[11] n17625_not ; n17626
g17371 and a[11] n17626_not ; n17627
g17372 and n17625_not n17626_not ; n17628
g17373 and n17627_not n17628_not ; n17629
g17374 and n17622_not n17629_not ; n17630
g17375 and n17622_not n17630_not ; n17631
g17376 and n17629_not n17630_not ; n17632
g17377 and n17631_not n17632_not ; n17633
g17378 and n17581_not n17585_not ; n17634
g17379 and b[62] n951 ; n17635
g17380 and b[60] n1056 ; n17636
g17381 and b[61] n946 ; n17637
g17382 and n17636_not n17637_not ; n17638
g17383 and n17635_not n17638 ; n17639
g17384 and n954_not n17639 ; n17640
g17385 and n13370_not n17639 ; n17641
g17386 and n17640_not n17641_not ; n17642
g17387 and a[14] n17642_not ; n17643
g17388 and a[14]_not n17642 ; n17644
g17389 and n17643_not n17644_not ; n17645
g17390 and n17634_not n17645_not ; n17646
g17391 and n17634 n17645 ; n17647
g17392 and n17646_not n17647_not ; n17648
g17393 and b[59] n1302 ; n17649
g17394 and b[57] n1391 ; n17650
g17395 and b[58] n1297 ; n17651
g17396 and n17650_not n17651_not ; n17652
g17397 and n17649_not n17652 ; n17653
g17398 and n1305 n12179 ; n17654
g17399 and n17653 n17654_not ; n17655
g17400 and a[17] n17655_not ; n17656
g17401 and a[17] n17656_not ; n17657
g17402 and n17655_not n17656_not ; n17658
g17403 and n17657_not n17658_not ; n17659
g17404 and n17287_not n17564_not ; n17660
g17405 and n17659 n17660 ; n17661
g17406 and n17659_not n17660_not ; n17662
g17407 and n17661_not n17662_not ; n17663
g17408 and b[56] n1627 ; n17664
g17409 and b[54] n1763 ; n17665
g17410 and b[55] n1622 ; n17666
g17411 and n17665_not n17666_not ; n17667
g17412 and n17664_not n17667 ; n17668
g17413 and n1630 n10708 ; n17669
g17414 and n17668 n17669_not ; n17670
g17415 and a[20] n17670_not ; n17671
g17416 and a[20] n17671_not ; n17672
g17417 and n17670_not n17671_not ; n17673
g17418 and n17672_not n17673_not ; n17674
g17419 and n17302_not n17561_not ; n17675
g17420 and n17674_not n17675_not ; n17676
g17421 and n17674_not n17676_not ; n17677
g17422 and n17675_not n17676_not ; n17678
g17423 and n17677_not n17678_not ; n17679
g17424 and n17549_not n17553_not ; n17680
g17425 and b[50] n2539 ; n17681
g17426 and b[48] n2685 ; n17682
g17427 and b[49] n2534 ; n17683
g17428 and n17682_not n17683_not ; n17684
g17429 and n17681_not n17684 ; n17685
g17430 and n2542_not n17685 ; n17686
g17431 and n8949_not n17685 ; n17687
g17432 and n17686_not n17687_not ; n17688
g17433 and a[26] n17688_not ; n17689
g17434 and a[26]_not n17688 ; n17690
g17435 and n17689_not n17690_not ; n17691
g17436 and n17680_not n17691_not ; n17692
g17437 and n17680 n17691 ; n17693
g17438 and n17692_not n17693_not ; n17694
g17439 and b[47] n3050 ; n17695
g17440 and b[45] n3243 ; n17696
g17441 and b[46] n3045 ; n17697
g17442 and n17696_not n17697_not ; n17698
g17443 and n17695_not n17698 ; n17699
g17444 and n3053 n7703 ; n17700
g17445 and n17699 n17700_not ; n17701
g17446 and a[29] n17701_not ; n17702
g17447 and a[29] n17702_not ; n17703
g17448 and n17701_not n17702_not ; n17704
g17449 and n17703_not n17704_not ; n17705
g17450 and n17334_not n17533_not ; n17706
g17451 and n17705 n17706 ; n17707
g17452 and n17705_not n17706_not ; n17708
g17453 and n17707_not n17708_not ; n17709
g17454 and n17525_not n17529_not ; n17710
g17455 and b[44] n3638 ; n17711
g17456 and b[42] n3843 ; n17712
g17457 and b[43] n3633 ; n17713
g17458 and n17712_not n17713_not ; n17714
g17459 and n17711_not n17714 ; n17715
g17460 and n3641_not n17715 ; n17716
g17461 and n7072_not n17715 ; n17717
g17462 and n17716_not n17717_not ; n17718
g17463 and a[32] n17718_not ; n17719
g17464 and a[32]_not n17718 ; n17720
g17465 and n17719_not n17720_not ; n17721
g17466 and n17710_not n17721_not ; n17722
g17467 and n17710 n17721 ; n17723
g17468 and n17722_not n17723_not ; n17724
g17469 and b[41] n4287 ; n17725
g17470 and b[39] n4532 ; n17726
g17471 and b[40] n4282 ; n17727
g17472 and n17726_not n17727_not ; n17728
g17473 and n17725_not n17728 ; n17729
g17474 and n4290 n6219 ; n17730
g17475 and n17729 n17730_not ; n17731
g17476 and a[35] n17731_not ; n17732
g17477 and a[35] n17732_not ; n17733
g17478 and n17731_not n17732_not ; n17734
g17479 and n17733_not n17734_not ; n17735
g17480 and n17517_not n17521_not ; n17736
g17481 and b[35] n5777 ; n17737
g17482 and b[33] n6059 ; n17738
g17483 and b[34] n5772 ; n17739
g17484 and n17738_not n17739_not ; n17740
g17485 and n17737_not n17740 ; n17741
g17486 and n4696 n5780 ; n17742
g17487 and n17741 n17742_not ; n17743
g17488 and a[41] n17743_not ; n17744
g17489 and a[41] n17744_not ; n17745
g17490 and n17743_not n17744_not ; n17746
g17491 and n17745_not n17746_not ; n17747
g17492 and n17457_not n17470_not ; n17748
g17493 and b[26] n8362 ; n17749
g17494 and b[24] n8715 ; n17750
g17495 and b[25] n8357 ; n17751
g17496 and n17750_not n17751_not ; n17752
g17497 and n17749_not n17752 ; n17753
g17498 and n2813 n8365 ; n17754
g17499 and n17753 n17754_not ; n17755
g17500 and a[50] n17755_not ; n17756
g17501 and a[50] n17756_not ; n17757
g17502 and n17755_not n17756_not ; n17758
g17503 and n17757_not n17758_not ; n17759
g17504 and n17438_not n17451_not ; n17760
g17505 and b[23] n9339 ; n17761
g17506 and b[21] n9732 ; n17762
g17507 and b[22] n9334 ; n17763
g17508 and n17762_not n17763_not ; n17764
g17509 and n17761_not n17764 ; n17765
g17510 and n2300 n9342 ; n17766
g17511 and n17765 n17766_not ; n17767
g17512 and a[53] n17767_not ; n17768
g17513 and a[53] n17768_not ; n17769
g17514 and n17767_not n17768_not ; n17770
g17515 and n17769_not n17770_not ; n17771
g17516 and n17419_not n17432_not ; n17772
g17517 and n17388_not n17392_not ; n17773
g17518 and b[10] n13903 ; n17774
g17519 and b[11] n13488_not ; n17775
g17520 and n17774_not n17775_not ; n17776
g17521 and n17385 n17776_not ; n17777
g17522 and n17385 n17777_not ; n17778
g17523 and n17776_not n17777_not ; n17779
g17524 and n17778_not n17779_not ; n17780
g17525 and n17773_not n17780_not ; n17781
g17526 and n17773_not n17781_not ; n17782
g17527 and n17780_not n17781_not ; n17783
g17528 and n17782_not n17783_not ; n17784
g17529 and b[14] n12668 ; n17785
g17530 and b[12] n13047 ; n17786
g17531 and b[13] n12663 ; n17787
g17532 and n17786_not n17787_not ; n17788
g17533 and n17785_not n17788 ; n17789
g17534 and n1034 n12671 ; n17790
g17535 and n17789 n17790_not ; n17791
g17536 and a[62] n17791_not ; n17792
g17537 and a[62] n17792_not ; n17793
g17538 and n17791_not n17792_not ; n17794
g17539 and n17793_not n17794_not ; n17795
g17540 and n17784_not n17795_not ; n17796
g17541 and n17784_not n17796_not ; n17797
g17542 and n17795_not n17796_not ; n17798
g17543 and n17797_not n17798_not ; n17799
g17544 and b[17] n11531 ; n17800
g17545 and b[15] n11896 ; n17801
g17546 and b[16] n11526 ; n17802
g17547 and n17801_not n17802_not ; n17803
g17548 and n17800_not n17803 ; n17804
g17549 and n1356 n11534 ; n17805
g17550 and n17804 n17805_not ; n17806
g17551 and a[59] n17806_not ; n17807
g17552 and a[59] n17807_not ; n17808
g17553 and n17806_not n17807_not ; n17809
g17554 and n17808_not n17809_not ; n17810
g17555 and n17799_not n17810_not ; n17811
g17556 and n17799_not n17811_not ; n17812
g17557 and n17810_not n17811_not ; n17813
g17558 and n17812_not n17813_not ; n17814
g17559 and n17398_not n17413_not ; n17815
g17560 and n17814 n17815 ; n17816
g17561 and n17814_not n17815_not ; n17817
g17562 and n17816_not n17817_not ; n17818
g17563 and b[20] n10426 ; n17819
g17564 and b[18] n10796 ; n17820
g17565 and b[19] n10421 ; n17821
g17566 and n17820_not n17821_not ; n17822
g17567 and n17819_not n17822 ; n17823
g17568 and n1846 n10429 ; n17824
g17569 and n17823 n17824_not ; n17825
g17570 and a[56] n17825_not ; n17826
g17571 and a[56] n17826_not ; n17827
g17572 and n17825_not n17826_not ; n17828
g17573 and n17827_not n17828_not ; n17829
g17574 and n17818_not n17829 ; n17830
g17575 and n17818 n17829_not ; n17831
g17576 and n17830_not n17831_not ; n17832
g17577 and n17772_not n17832 ; n17833
g17578 and n17772_not n17833_not ; n17834
g17579 and n17832 n17833_not ; n17835
g17580 and n17834_not n17835_not ; n17836
g17581 and n17771_not n17836_not ; n17837
g17582 and n17771 n17835_not ; n17838
g17583 and n17834_not n17838 ; n17839
g17584 and n17837_not n17839_not ; n17840
g17585 and n17760_not n17840 ; n17841
g17586 and n17760 n17840_not ; n17842
g17587 and n17841_not n17842_not ; n17843
g17588 and n17759_not n17843 ; n17844
g17589 and n17759 n17843_not ; n17845
g17590 and n17844_not n17845_not ; n17846
g17591 and n17748_not n17846 ; n17847
g17592 and n17748 n17846_not ; n17848
g17593 and n17847_not n17848_not ; n17849
g17594 and b[29] n7446 ; n17850
g17595 and b[27] n7787 ; n17851
g17596 and b[28] n7441 ; n17852
g17597 and n17851_not n17852_not ; n17853
g17598 and n17850_not n17853 ; n17854
g17599 and n3383 n7449 ; n17855
g17600 and n17854 n17855_not ; n17856
g17601 and a[47] n17856_not ; n17857
g17602 and a[47] n17857_not ; n17858
g17603 and n17856_not n17857_not ; n17859
g17604 and n17858_not n17859_not ; n17860
g17605 and n17849 n17860_not ; n17861
g17606 and n17849 n17861_not ; n17862
g17607 and n17860_not n17861_not ; n17863
g17608 and n17862_not n17863_not ; n17864
g17609 and n17476_not n17489_not ; n17865
g17610 and n17864 n17865 ; n17866
g17611 and n17864_not n17865_not ; n17867
g17612 and n17866_not n17867_not ; n17868
g17613 and b[32] n6595 ; n17869
g17614 and b[30] n6902 ; n17870
g17615 and b[31] n6590 ; n17871
g17616 and n17870_not n17871_not ; n17872
g17617 and n17869_not n17872 ; n17873
g17618 and n4013 n6598 ; n17874
g17619 and n17873 n17874_not ; n17875
g17620 and a[44] n17875_not ; n17876
g17621 and a[44] n17876_not ; n17877
g17622 and n17875_not n17876_not ; n17878
g17623 and n17877_not n17878_not ; n17879
g17624 and n17868_not n17879 ; n17880
g17625 and n17868 n17879_not ; n17881
g17626 and n17880_not n17881_not ; n17882
g17627 and n17495_not n17509_not ; n17883
g17628 and n17882 n17883_not ; n17884
g17629 and n17882_not n17883 ; n17885
g17630 and n17884_not n17885_not ; n17886
g17631 and n17747_not n17886 ; n17887
g17632 and n17886 n17887_not ; n17888
g17633 and n17747_not n17887_not ; n17889
g17634 and n17888_not n17889_not ; n17890
g17635 and n17511_not n17514_not ; n17891
g17636 and n17890 n17891 ; n17892
g17637 and n17890_not n17891_not ; n17893
g17638 and n17892_not n17893_not ; n17894
g17639 and b[38] n5035 ; n17895
g17640 and b[36] n5277 ; n17896
g17641 and b[37] n5030 ; n17897
g17642 and n17896_not n17897_not ; n17898
g17643 and n17895_not n17898 ; n17899
g17644 and n5038 n5205 ; n17900
g17645 and n17899 n17900_not ; n17901
g17646 and a[38] n17901_not ; n17902
g17647 and a[38] n17902_not ; n17903
g17648 and n17901_not n17902_not ; n17904
g17649 and n17903_not n17904_not ; n17905
g17650 and n17894_not n17905 ; n17906
g17651 and n17894 n17905_not ; n17907
g17652 and n17906_not n17907_not ; n17908
g17653 and n17736_not n17908 ; n17909
g17654 and n17736 n17908_not ; n17910
g17655 and n17909_not n17910_not ; n17911
g17656 and n17735_not n17911 ; n17912
g17657 and n17735_not n17912_not ; n17913
g17658 and n17911 n17912_not ; n17914
g17659 and n17913_not n17914_not ; n17915
g17660 and n17724 n17915_not ; n17916
g17661 and n17724 n17916_not ; n17917
g17662 and n17915_not n17916_not ; n17918
g17663 and n17917_not n17918_not ; n17919
g17664 and n17709 n17919_not ; n17920
g17665 and n17709_not n17919 ; n17921
g17666 and n17694 n17921_not ; n17922
g17667 and n17920_not n17922 ; n17923
g17668 and n17694 n17923_not ; n17924
g17669 and n17921_not n17923_not ; n17925
g17670 and n17920_not n17925 ; n17926
g17671 and n17924_not n17926_not ; n17927
g17672 and n17317_not n17557_not ; n17928
g17673 and b[53] n2048 ; n17929
g17674 and b[51] n2198 ; n17930
g17675 and b[52] n2043 ; n17931
g17676 and n17930_not n17931_not ; n17932
g17677 and n17929_not n17932 ; n17933
g17678 and n2051_not n17933 ; n17934
g17679 and n9972_not n17933 ; n17935
g17680 and n17934_not n17935_not ; n17936
g17681 and a[23] n17936_not ; n17937
g17682 and a[23]_not n17936 ; n17938
g17683 and n17937_not n17938_not ; n17939
g17684 and n17928_not n17939_not ; n17940
g17685 and n17928_not n17940_not ; n17941
g17686 and n17939_not n17940_not ; n17942
g17687 and n17941_not n17942_not ; n17943
g17688 and n17927_not n17943_not ; n17944
g17689 and n17927_not n17944_not ; n17945
g17690 and n17943_not n17944_not ; n17946
g17691 and n17945_not n17946_not ; n17947
g17692 and n17679_not n17947_not ; n17948
g17693 and n17679_not n17948_not ; n17949
g17694 and n17947_not n17948_not ; n17950
g17695 and n17949_not n17950_not ; n17951
g17696 and n17663 n17951_not ; n17952
g17697 and n17663_not n17951 ; n17953
g17698 and n17648 n17953_not ; n17954
g17699 and n17952_not n17954 ; n17955
g17700 and n17648 n17955_not ; n17956
g17701 and n17953_not n17955_not ; n17957
g17702 and n17952_not n17957 ; n17958
g17703 and n17956_not n17958_not ; n17959
g17704 and n17633_not n17959 ; n17960
g17705 and n17633 n17959_not ; n17961
g17706 and n17960_not n17961_not ; n17962
g17707 and n17621_not n17962_not ; n17963
g17708 and n17621_not n17963_not ; n17964
g17709 and n17962_not n17963_not ; n17965
g17710 and n17964_not n17965_not ; n17966
g17711 and n17620_not n17966_not ; n17967
g17712 and n17620 n17965_not ; n17968
g17713 and n17964_not n17968 ; n17969
g17714 and n17967_not n17969_not ; f[74]
g17715 and n17963_not n17967_not ; n17971
g17716 and n17633_not n17959_not ; n17972
g17717 and n17630_not n17972_not ; n17973
g17718 and n17646_not n17955_not ; n17974
g17719 and b[63] n951 ; n17975
g17720 and b[61] n1056 ; n17976
g17721 and b[62] n946 ; n17977
g17722 and n17976_not n17977_not ; n17978
g17723 and n17975_not n17978 ; n17979
g17724 and n954 n13771 ; n17980
g17725 and n17979 n17980_not ; n17981
g17726 and a[14] n17981_not ; n17982
g17727 and a[14] n17982_not ; n17983
g17728 and n17981_not n17982_not ; n17984
g17729 and n17983_not n17984_not ; n17985
g17730 and n17974_not n17985_not ; n17986
g17731 and n17974_not n17986_not ; n17987
g17732 and n17985_not n17986_not ; n17988
g17733 and n17987_not n17988_not ; n17989
g17734 and n17662_not n17952_not ; n17990
g17735 and b[60] n1302 ; n17991
g17736 and b[58] n1391 ; n17992
g17737 and b[59] n1297 ; n17993
g17738 and n17992_not n17993_not ; n17994
g17739 and n17991_not n17994 ; n17995
g17740 and n1305 n12211 ; n17996
g17741 and n17995 n17996_not ; n17997
g17742 and a[17] n17997_not ; n17998
g17743 and a[17] n17998_not ; n17999
g17744 and n17997_not n17998_not ; n18000
g17745 and n17999_not n18000_not ; n18001
g17746 and n17990_not n18001 ; n18002
g17747 and n17990 n18001_not ; n18003
g17748 and n18002_not n18003_not ; n18004
g17749 and b[57] n1627 ; n18005
g17750 and b[55] n1763 ; n18006
g17751 and b[56] n1622 ; n18007
g17752 and n18006_not n18007_not ; n18008
g17753 and n18005_not n18008 ; n18009
g17754 and n1630 n11410 ; n18010
g17755 and n18009 n18010_not ; n18011
g17756 and a[20] n18011_not ; n18012
g17757 and a[20] n18012_not ; n18013
g17758 and n18011_not n18012_not ; n18014
g17759 and n18013_not n18014_not ; n18015
g17760 and n17676_not n17948_not ; n18016
g17761 and n18015 n18016 ; n18017
g17762 and n18015_not n18016_not ; n18018
g17763 and n18017_not n18018_not ; n18019
g17764 and n17940_not n17944_not ; n18020
g17765 and b[54] n2048 ; n18021
g17766 and b[52] n2198 ; n18022
g17767 and b[53] n2043 ; n18023
g17768 and n18022_not n18023_not ; n18024
g17769 and n18021_not n18024 ; n18025
g17770 and n2051 n9998 ; n18026
g17771 and n18025 n18026_not ; n18027
g17772 and a[23] n18027_not ; n18028
g17773 and a[23] n18028_not ; n18029
g17774 and n18027_not n18028_not ; n18030
g17775 and n18029_not n18030_not ; n18031
g17776 and n18020_not n18031_not ; n18032
g17777 and n18020_not n18032_not ; n18033
g17778 and n18031_not n18032_not ; n18034
g17779 and n18033_not n18034_not ; n18035
g17780 and b[51] n2539 ; n18036
g17781 and b[49] n2685 ; n18037
g17782 and b[50] n2534 ; n18038
g17783 and n18037_not n18038_not ; n18039
g17784 and n18036_not n18039 ; n18040
g17785 and n2542 n8976 ; n18041
g17786 and n18040 n18041_not ; n18042
g17787 and a[26] n18042_not ; n18043
g17788 and a[26] n18043_not ; n18044
g17789 and n18042_not n18043_not ; n18045
g17790 and n18044_not n18045_not ; n18046
g17791 and n17692_not n17923_not ; n18047
g17792 and n18046 n18047 ; n18048
g17793 and n18046_not n18047_not ; n18049
g17794 and n18048_not n18049_not ; n18050
g17795 and n17708_not n17920_not ; n18051
g17796 and b[48] n3050 ; n18052
g17797 and b[46] n3243 ; n18053
g17798 and b[47] n3045 ; n18054
g17799 and n18053_not n18054_not ; n18055
g17800 and n18052_not n18055 ; n18056
g17801 and n3053 n8009 ; n18057
g17802 and n18056 n18057_not ; n18058
g17803 and a[29] n18058_not ; n18059
g17804 and a[29] n18059_not ; n18060
g17805 and n18058_not n18059_not ; n18061
g17806 and n18060_not n18061_not ; n18062
g17807 and n18051_not n18062 ; n18063
g17808 and n18051 n18062_not ; n18064
g17809 and n18063_not n18064_not ; n18065
g17810 and n17909_not n17912_not ; n18066
g17811 and n17893_not n17907_not ; n18067
g17812 and n17884_not n17887_not ; n18068
g17813 and n17867_not n17881_not ; n18069
g17814 and n17847_not n17861_not ; n18070
g17815 and n17833_not n17837_not ; n18071
g17816 and b[24] n9339 ; n18072
g17817 and b[22] n9732 ; n18073
g17818 and b[23] n9334 ; n18074
g17819 and n18073_not n18074_not ; n18075
g17820 and n18072_not n18075 ; n18076
g17821 and n2458 n9342 ; n18077
g17822 and n18076 n18077_not ; n18078
g17823 and a[53] n18078_not ; n18079
g17824 and a[53] n18079_not ; n18080
g17825 and n18078_not n18079_not ; n18081
g17826 and n18080_not n18081_not ; n18082
g17827 and n17777_not n17781_not ; n18083
g17828 and b[15] n12668 ; n18084
g17829 and b[13] n13047 ; n18085
g17830 and b[14] n12663 ; n18086
g17831 and n18085_not n18086_not ; n18087
g17832 and n18084_not n18087 ; n18088
g17833 and n1131 n12671 ; n18089
g17834 and n18088 n18089_not ; n18090
g17835 and a[62] n18090_not ; n18091
g17836 and a[62] n18091_not ; n18092
g17837 and n18090_not n18091_not ; n18093
g17838 and n18092_not n18093_not ; n18094
g17839 and b[11] n13903 ; n18095
g17840 and b[12] n13488_not ; n18096
g17841 and n18095_not n18096_not ; n18097
g17842 and a[11] n17385_not ; n18098
g17843 and a[11]_not n17385 ; n18099
g17844 and n18098_not n18099_not ; n18100
g17845 and n18097_not n18100_not ; n18101
g17846 and n18097 n18100 ; n18102
g17847 and n18101_not n18102_not ; n18103
g17848 and n18094_not n18103 ; n18104
g17849 and n18094_not n18104_not ; n18105
g17850 and n18103 n18104_not ; n18106
g17851 and n18105_not n18106_not ; n18107
g17852 and n18083_not n18107_not ; n18108
g17853 and n18083_not n18108_not ; n18109
g17854 and n18107_not n18108_not ; n18110
g17855 and n18109_not n18110_not ; n18111
g17856 and b[18] n11531 ; n18112
g17857 and b[16] n11896 ; n18113
g17858 and b[17] n11526 ; n18114
g17859 and n18113_not n18114_not ; n18115
g17860 and n18112_not n18115 ; n18116
g17861 and n1566 n11534 ; n18117
g17862 and n18116 n18117_not ; n18118
g17863 and a[59] n18118_not ; n18119
g17864 and a[59] n18119_not ; n18120
g17865 and n18118_not n18119_not ; n18121
g17866 and n18120_not n18121_not ; n18122
g17867 and n18111_not n18122_not ; n18123
g17868 and n18111_not n18123_not ; n18124
g17869 and n18122_not n18123_not ; n18125
g17870 and n18124_not n18125_not ; n18126
g17871 and n17796_not n17811_not ; n18127
g17872 and n18126 n18127 ; n18128
g17873 and n18126_not n18127_not ; n18129
g17874 and n18128_not n18129_not ; n18130
g17875 and b[21] n10426 ; n18131
g17876 and b[19] n10796 ; n18132
g17877 and b[20] n10421 ; n18133
g17878 and n18132_not n18133_not ; n18134
g17879 and n18131_not n18134 ; n18135
g17880 and n1984 n10429 ; n18136
g17881 and n18135 n18136_not ; n18137
g17882 and a[56] n18137_not ; n18138
g17883 and a[56] n18138_not ; n18139
g17884 and n18137_not n18138_not ; n18140
g17885 and n18139_not n18140_not ; n18141
g17886 and n18130 n18141_not ; n18142
g17887 and n18130 n18142_not ; n18143
g17888 and n18141_not n18142_not ; n18144
g17889 and n18143_not n18144_not ; n18145
g17890 and n17817_not n17831_not ; n18146
g17891 and n18145_not n18146_not ; n18147
g17892 and n18145 n18146 ; n18148
g17893 and n18147_not n18148_not ; n18149
g17894 and n18082_not n18149 ; n18150
g17895 and n18082_not n18150_not ; n18151
g17896 and n18149 n18150_not ; n18152
g17897 and n18151_not n18152_not ; n18153
g17898 and n18071_not n18153_not ; n18154
g17899 and n18071_not n18154_not ; n18155
g17900 and n18153_not n18154_not ; n18156
g17901 and n18155_not n18156_not ; n18157
g17902 and b[27] n8362 ; n18158
g17903 and b[25] n8715 ; n18159
g17904 and b[26] n8357 ; n18160
g17905 and n18159_not n18160_not ; n18161
g17906 and n18158_not n18161 ; n18162
g17907 and n2990 n8365 ; n18163
g17908 and n18162 n18163_not ; n18164
g17909 and a[50] n18164_not ; n18165
g17910 and a[50] n18165_not ; n18166
g17911 and n18164_not n18165_not ; n18167
g17912 and n18166_not n18167_not ; n18168
g17913 and n18157_not n18168_not ; n18169
g17914 and n18157_not n18169_not ; n18170
g17915 and n18168_not n18169_not ; n18171
g17916 and n18170_not n18171_not ; n18172
g17917 and n17841_not n17844_not ; n18173
g17918 and n18172 n18173 ; n18174
g17919 and n18172_not n18173_not ; n18175
g17920 and n18174_not n18175_not ; n18176
g17921 and b[30] n7446 ; n18177
g17922 and b[28] n7787 ; n18178
g17923 and b[29] n7441 ; n18179
g17924 and n18178_not n18179_not ; n18180
g17925 and n18177_not n18180 ; n18181
g17926 and n3577 n7449 ; n18182
g17927 and n18181 n18182_not ; n18183
g17928 and a[47] n18183_not ; n18184
g17929 and a[47] n18184_not ; n18185
g17930 and n18183_not n18184_not ; n18186
g17931 and n18185_not n18186_not ; n18187
g17932 and n18176 n18187_not ; n18188
g17933 and n18176_not n18187 ; n18189
g17934 and n18070_not n18189_not ; n18190
g17935 and n18188_not n18190 ; n18191
g17936 and n18070_not n18191_not ; n18192
g17937 and n18188_not n18191_not ; n18193
g17938 and n18189_not n18193 ; n18194
g17939 and n18192_not n18194_not ; n18195
g17940 and b[33] n6595 ; n18196
g17941 and b[31] n6902 ; n18197
g17942 and b[32] n6590 ; n18198
g17943 and n18197_not n18198_not ; n18199
g17944 and n18196_not n18199 ; n18200
g17945 and n4223 n6598 ; n18201
g17946 and n18200 n18201_not ; n18202
g17947 and a[44] n18202_not ; n18203
g17948 and a[44] n18203_not ; n18204
g17949 and n18202_not n18203_not ; n18205
g17950 and n18204_not n18205_not ; n18206
g17951 and n18195_not n18206_not ; n18207
g17952 and n18195_not n18207_not ; n18208
g17953 and n18206_not n18207_not ; n18209
g17954 and n18208_not n18209_not ; n18210
g17955 and n18069_not n18210 ; n18211
g17956 and n18069 n18210_not ; n18212
g17957 and n18211_not n18212_not ; n18213
g17958 and b[36] n5777 ; n18214
g17959 and b[34] n6059 ; n18215
g17960 and b[35] n5772 ; n18216
g17961 and n18215_not n18216_not ; n18217
g17962 and n18214_not n18217 ; n18218
g17963 and n4922 n5780 ; n18219
g17964 and n18218 n18219_not ; n18220
g17965 and a[41] n18220_not ; n18221
g17966 and a[41] n18221_not ; n18222
g17967 and n18220_not n18221_not ; n18223
g17968 and n18222_not n18223_not ; n18224
g17969 and n18213_not n18224_not ; n18225
g17970 and n18213 n18224 ; n18226
g17971 and n18225_not n18226_not ; n18227
g17972 and n18068 n18227_not ; n18228
g17973 and n18068_not n18227 ; n18229
g17974 and n18228_not n18229_not ; n18230
g17975 and b[39] n5035 ; n18231
g17976 and b[37] n5277 ; n18232
g17977 and b[38] n5030 ; n18233
g17978 and n18232_not n18233_not ; n18234
g17979 and n18231_not n18234 ; n18235
g17980 and n5038 n5451 ; n18236
g17981 and n18235 n18236_not ; n18237
g17982 and a[38] n18237_not ; n18238
g17983 and a[38] n18238_not ; n18239
g17984 and n18237_not n18238_not ; n18240
g17985 and n18239_not n18240_not ; n18241
g17986 and n18230 n18241_not ; n18242
g17987 and n18230 n18242_not ; n18243
g17988 and n18241_not n18242_not ; n18244
g17989 and n18243_not n18244_not ; n18245
g17990 and n18067_not n18245 ; n18246
g17991 and n18067 n18245_not ; n18247
g17992 and n18246_not n18247_not ; n18248
g17993 and b[42] n4287 ; n18249
g17994 and b[40] n4532 ; n18250
g17995 and b[41] n4282 ; n18251
g17996 and n18250_not n18251_not ; n18252
g17997 and n18249_not n18252 ; n18253
g17998 and n4290 n6489 ; n18254
g17999 and n18253 n18254_not ; n18255
g18000 and a[35] n18255_not ; n18256
g18001 and a[35] n18256_not ; n18257
g18002 and n18255_not n18256_not ; n18258
g18003 and n18257_not n18258_not ; n18259
g18004 and n18248_not n18259_not ; n18260
g18005 and n18248 n18259 ; n18261
g18006 and n18260_not n18261_not ; n18262
g18007 and n18066 n18262_not ; n18263
g18008 and n18066_not n18262 ; n18264
g18009 and n18263_not n18264_not ; n18265
g18010 and n17722_not n17916_not ; n18266
g18011 and b[45] n3638 ; n18267
g18012 and b[43] n3843 ; n18268
g18013 and b[44] n3633 ; n18269
g18014 and n18268_not n18269_not ; n18270
g18015 and n18267_not n18270 ; n18271
g18016 and n3641 n7361 ; n18272
g18017 and n18271 n18272_not ; n18273
g18018 and a[32] n18273_not ; n18274
g18019 and a[32] n18274_not ; n18275
g18020 and n18273_not n18274_not ; n18276
g18021 and n18275_not n18276_not ; n18277
g18022 and n18266_not n18277_not ; n18278
g18023 and n18266_not n18278_not ; n18279
g18024 and n18277_not n18278_not ; n18280
g18025 and n18279_not n18280_not ; n18281
g18026 and n18265 n18281_not ; n18282
g18027 and n18265_not n18281 ; n18283
g18028 and n18065_not n18283_not ; n18284
g18029 and n18282_not n18284 ; n18285
g18030 and n18065_not n18285_not ; n18286
g18031 and n18283_not n18285_not ; n18287
g18032 and n18282_not n18287 ; n18288
g18033 and n18286_not n18288_not ; n18289
g18034 and n18050 n18289_not ; n18290
g18035 and n18050_not n18289 ; n18291
g18036 and n18035_not n18291_not ; n18292
g18037 and n18290_not n18292 ; n18293
g18038 and n18035_not n18293_not ; n18294
g18039 and n18291_not n18293_not ; n18295
g18040 and n18290_not n18295 ; n18296
g18041 and n18294_not n18296_not ; n18297
g18042 and n18019 n18297_not ; n18298
g18043 and n18019_not n18297 ; n18299
g18044 and n18004_not n18299_not ; n18300
g18045 and n18298_not n18300 ; n18301
g18046 and n18004_not n18301_not ; n18302
g18047 and n18299_not n18301_not ; n18303
g18048 and n18298_not n18303 ; n18304
g18049 and n18302_not n18304_not ; n18305
g18050 and n17989_not n18305 ; n18306
g18051 and n17989 n18305_not ; n18307
g18052 and n18306_not n18307_not ; n18308
g18053 and n17973_not n18308_not ; n18309
g18054 and n17973_not n18309_not ; n18310
g18055 and n18308_not n18309_not ; n18311
g18056 and n18310_not n18311_not ; n18312
g18057 and n17971_not n18312_not ; n18313
g18058 and n17971 n18311_not ; n18314
g18059 and n18310_not n18314 ; n18315
g18060 and n18313_not n18315_not ; f[75]
g18061 and n18309_not n18313_not ; n18317
g18062 and n17989_not n18305_not ; n18318
g18063 and n17986_not n18318_not ; n18319
g18064 and b[61] n1302 ; n18320
g18065 and b[59] n1391 ; n18321
g18066 and b[60] n1297 ; n18322
g18067 and n18321_not n18322_not ; n18323
g18068 and n18320_not n18323 ; n18324
g18069 and n1305 n12969 ; n18325
g18070 and n18324 n18325_not ; n18326
g18071 and a[17] n18326_not ; n18327
g18072 and a[17] n18327_not ; n18328
g18073 and n18326_not n18327_not ; n18329
g18074 and n18328_not n18329_not ; n18330
g18075 and n18018_not n18298_not ; n18331
g18076 and n18330_not n18331_not ; n18332
g18077 and n18330_not n18332_not ; n18333
g18078 and n18331_not n18332_not ; n18334
g18079 and n18333_not n18334_not ; n18335
g18080 and b[55] n2048 ; n18336
g18081 and b[53] n2198 ; n18337
g18082 and b[54] n2043 ; n18338
g18083 and n18337_not n18338_not ; n18339
g18084 and n18336_not n18339 ; n18340
g18085 and n2051 n10684 ; n18341
g18086 and n18340 n18341_not ; n18342
g18087 and a[23] n18342_not ; n18343
g18088 and a[23] n18343_not ; n18344
g18089 and n18342_not n18343_not ; n18345
g18090 and n18344_not n18345_not ; n18346
g18091 and n18049_not n18290_not ; n18347
g18092 and n18346_not n18347_not ; n18348
g18093 and n18346_not n18348_not ; n18349
g18094 and n18347_not n18348_not ; n18350
g18095 and n18349_not n18350_not ; n18351
g18096 and b[49] n3050 ; n18352
g18097 and b[47] n3243 ; n18353
g18098 and b[48] n3045 ; n18354
g18099 and n18353_not n18354_not ; n18355
g18100 and n18352_not n18355 ; n18356
g18101 and n3053 n8625 ; n18357
g18102 and n18356 n18357_not ; n18358
g18103 and a[29] n18358_not ; n18359
g18104 and a[29] n18359_not ; n18360
g18105 and n18358_not n18359_not ; n18361
g18106 and n18360_not n18361_not ; n18362
g18107 and n18278_not n18282_not ; n18363
g18108 and n18362_not n18363_not ; n18364
g18109 and n18362_not n18364_not ; n18365
g18110 and n18363_not n18364_not ; n18366
g18111 and n18365_not n18366_not ; n18367
g18112 and b[43] n4287 ; n18368
g18113 and b[41] n4532 ; n18369
g18114 and b[42] n4282 ; n18370
g18115 and n18369_not n18370_not ; n18371
g18116 and n18368_not n18371 ; n18372
g18117 and n4290 n6515 ; n18373
g18118 and n18372 n18373_not ; n18374
g18119 and a[35] n18374_not ; n18375
g18120 and a[35] n18375_not ; n18376
g18121 and n18374_not n18375_not ; n18377
g18122 and n18376_not n18377_not ; n18378
g18123 and n18067_not n18245_not ; n18379
g18124 and n18242_not n18379_not ; n18380
g18125 and b[40] n5035 ; n18381
g18126 and b[38] n5277 ; n18382
g18127 and b[39] n5030 ; n18383
g18128 and n18382_not n18383_not ; n18384
g18129 and n18381_not n18384 ; n18385
g18130 and n5038 n5955 ; n18386
g18131 and n18385 n18386_not ; n18387
g18132 and a[38] n18387_not ; n18388
g18133 and a[38] n18388_not ; n18389
g18134 and n18387_not n18388_not ; n18390
g18135 and n18389_not n18390_not ; n18391
g18136 and n18225_not n18229_not ; n18392
g18137 and b[37] n5777 ; n18393
g18138 and b[35] n6059 ; n18394
g18139 and b[36] n5772 ; n18395
g18140 and n18394_not n18395_not ; n18396
g18141 and n18393_not n18396 ; n18397
g18142 and n5181 n5780 ; n18398
g18143 and n18397 n18398_not ; n18399
g18144 and a[41] n18399_not ; n18400
g18145 and a[41] n18400_not ; n18401
g18146 and n18399_not n18400_not ; n18402
g18147 and n18401_not n18402_not ; n18403
g18148 and n18069_not n18210_not ; n18404
g18149 and n18207_not n18404_not ; n18405
g18150 and b[34] n6595 ; n18406
g18151 and b[32] n6902 ; n18407
g18152 and b[33] n6590 ; n18408
g18153 and n18407_not n18408_not ; n18409
g18154 and n18406_not n18409 ; n18410
g18155 and n4466 n6598 ; n18411
g18156 and n18410 n18411_not ; n18412
g18157 and a[44] n18412_not ; n18413
g18158 and a[44] n18413_not ; n18414
g18159 and n18412_not n18413_not ; n18415
g18160 and n18414_not n18415_not ; n18416
g18161 and b[31] n7446 ; n18417
g18162 and b[29] n7787 ; n18418
g18163 and b[30] n7441 ; n18419
g18164 and n18418_not n18419_not ; n18420
g18165 and n18417_not n18420 ; n18421
g18166 and n3796 n7449 ; n18422
g18167 and n18421 n18422_not ; n18423
g18168 and a[47] n18423_not ; n18424
g18169 and a[47] n18424_not ; n18425
g18170 and n18423_not n18424_not ; n18426
g18171 and n18425_not n18426_not ; n18427
g18172 and n18169_not n18175_not ; n18428
g18173 and b[12] n13903 ; n18429
g18174 and b[13] n13488_not ; n18430
g18175 and n18429_not n18430_not ; n18431
g18176 and a[11]_not n17385_not ; n18432
g18177 and n18101_not n18432_not ; n18433
g18178 and n18431 n18433_not ; n18434
g18179 and n18431 n18434_not ; n18435
g18180 and n18433_not n18434_not ; n18436
g18181 and n18435_not n18436_not ; n18437
g18182 and b[16] n12668 ; n18438
g18183 and b[14] n13047 ; n18439
g18184 and b[15] n12663 ; n18440
g18185 and n18439_not n18440_not ; n18441
g18186 and n18438_not n18441 ; n18442
g18187 and n1237 n12671 ; n18443
g18188 and n18442 n18443_not ; n18444
g18189 and a[62] n18444_not ; n18445
g18190 and a[62] n18445_not ; n18446
g18191 and n18444_not n18445_not ; n18447
g18192 and n18446_not n18447_not ; n18448
g18193 and n18437_not n18448 ; n18449
g18194 and n18437 n18448_not ; n18450
g18195 and n18449_not n18450_not ; n18451
g18196 and n18104_not n18108_not ; n18452
g18197 and n18451 n18452 ; n18453
g18198 and n18451_not n18452_not ; n18454
g18199 and n18453_not n18454_not ; n18455
g18200 and b[19] n11531 ; n18456
g18201 and b[17] n11896 ; n18457
g18202 and b[18] n11526 ; n18458
g18203 and n18457_not n18458_not ; n18459
g18204 and n18456_not n18459 ; n18460
g18205 and n1708 n11534 ; n18461
g18206 and n18460 n18461_not ; n18462
g18207 and a[59] n18462_not ; n18463
g18208 and a[59] n18463_not ; n18464
g18209 and n18462_not n18463_not ; n18465
g18210 and n18464_not n18465_not ; n18466
g18211 and n18455 n18466_not ; n18467
g18212 and n18455 n18467_not ; n18468
g18213 and n18466_not n18467_not ; n18469
g18214 and n18468_not n18469_not ; n18470
g18215 and n18123_not n18129_not ; n18471
g18216 and n18470 n18471 ; n18472
g18217 and n18470_not n18471_not ; n18473
g18218 and n18472_not n18473_not ; n18474
g18219 and b[22] n10426 ; n18475
g18220 and b[20] n10796 ; n18476
g18221 and b[21] n10421 ; n18477
g18222 and n18476_not n18477_not ; n18478
g18223 and n18475_not n18478 ; n18479
g18224 and n2145 n10429 ; n18480
g18225 and n18479 n18480_not ; n18481
g18226 and a[56] n18481_not ; n18482
g18227 and a[56] n18482_not ; n18483
g18228 and n18481_not n18482_not ; n18484
g18229 and n18483_not n18484_not ; n18485
g18230 and n18474 n18485_not ; n18486
g18231 and n18474 n18486_not ; n18487
g18232 and n18485_not n18486_not ; n18488
g18233 and n18487_not n18488_not ; n18489
g18234 and n18142_not n18147_not ; n18490
g18235 and n18489 n18490 ; n18491
g18236 and n18489_not n18490_not ; n18492
g18237 and n18491_not n18492_not ; n18493
g18238 and b[25] n9339 ; n18494
g18239 and b[23] n9732 ; n18495
g18240 and b[24] n9334 ; n18496
g18241 and n18495_not n18496_not ; n18497
g18242 and n18494_not n18497 ; n18498
g18243 and n2485 n9342 ; n18499
g18244 and n18498 n18499_not ; n18500
g18245 and a[53] n18500_not ; n18501
g18246 and a[53] n18501_not ; n18502
g18247 and n18500_not n18501_not ; n18503
g18248 and n18502_not n18503_not ; n18504
g18249 and n18493 n18504_not ; n18505
g18250 and n18493 n18505_not ; n18506
g18251 and n18504_not n18505_not ; n18507
g18252 and n18506_not n18507_not ; n18508
g18253 and n18150_not n18154_not ; n18509
g18254 and n18508 n18509 ; n18510
g18255 and n18508_not n18509_not ; n18511
g18256 and n18510_not n18511_not ; n18512
g18257 and b[28] n8362 ; n18513
g18258 and b[26] n8715 ; n18514
g18259 and b[27] n8357 ; n18515
g18260 and n18514_not n18515_not ; n18516
g18261 and n18513_not n18516 ; n18517
g18262 and n3189 n8365 ; n18518
g18263 and n18517 n18518_not ; n18519
g18264 and a[50] n18519_not ; n18520
g18265 and a[50] n18520_not ; n18521
g18266 and n18519_not n18520_not ; n18522
g18267 and n18521_not n18522_not ; n18523
g18268 and n18512_not n18523 ; n18524
g18269 and n18512 n18523_not ; n18525
g18270 and n18524_not n18525_not ; n18526
g18271 and n18428_not n18526 ; n18527
g18272 and n18428_not n18527_not ; n18528
g18273 and n18526 n18527_not ; n18529
g18274 and n18528_not n18529_not ; n18530
g18275 and n18427_not n18530_not ; n18531
g18276 and n18427 n18529_not ; n18532
g18277 and n18528_not n18532 ; n18533
g18278 and n18531_not n18533_not ; n18534
g18279 and n18193_not n18534 ; n18535
g18280 and n18193 n18534_not ; n18536
g18281 and n18535_not n18536_not ; n18537
g18282 and n18416_not n18537 ; n18538
g18283 and n18416 n18537_not ; n18539
g18284 and n18538_not n18539_not ; n18540
g18285 and n18405_not n18540 ; n18541
g18286 and n18405_not n18541_not ; n18542
g18287 and n18540 n18541_not ; n18543
g18288 and n18542_not n18543_not ; n18544
g18289 and n18403_not n18544_not ; n18545
g18290 and n18403 n18543_not ; n18546
g18291 and n18542_not n18546 ; n18547
g18292 and n18545_not n18547_not ; n18548
g18293 and n18392_not n18548 ; n18549
g18294 and n18392_not n18549_not ; n18550
g18295 and n18548 n18549_not ; n18551
g18296 and n18550_not n18551_not ; n18552
g18297 and n18391_not n18552_not ; n18553
g18298 and n18391 n18551_not ; n18554
g18299 and n18550_not n18554 ; n18555
g18300 and n18553_not n18555_not ; n18556
g18301 and n18380_not n18556 ; n18557
g18302 and n18380 n18556_not ; n18558
g18303 and n18557_not n18558_not ; n18559
g18304 and n18378_not n18559 ; n18560
g18305 and n18559 n18560_not ; n18561
g18306 and n18378_not n18560_not ; n18562
g18307 and n18561_not n18562_not ; n18563
g18308 and n18260_not n18264_not ; n18564
g18309 and b[46] n3638 ; n18565
g18310 and b[44] n3843 ; n18566
g18311 and b[45] n3633 ; n18567
g18312 and n18566_not n18567_not ; n18568
g18313 and n18565_not n18568 ; n18569
g18314 and n3641_not n18569 ; n18570
g18315 and n7677_not n18569 ; n18571
g18316 and n18570_not n18571_not ; n18572
g18317 and a[32] n18572_not ; n18573
g18318 and a[32]_not n18572 ; n18574
g18319 and n18573_not n18574_not ; n18575
g18320 and n18564_not n18575_not ; n18576
g18321 and n18564_not n18576_not ; n18577
g18322 and n18575_not n18576_not ; n18578
g18323 and n18577_not n18578_not ; n18579
g18324 and n18563_not n18579_not ; n18580
g18325 and n18563_not n18580_not ; n18581
g18326 and n18579_not n18580_not ; n18582
g18327 and n18581_not n18582_not ; n18583
g18328 and n18367_not n18583_not ; n18584
g18329 and n18367_not n18584_not ; n18585
g18330 and n18583_not n18584_not ; n18586
g18331 and n18585_not n18586_not ; n18587
g18332 and n18051_not n18062_not ; n18588
g18333 and n18285_not n18588_not ; n18589
g18334 and b[52] n2539 ; n18590
g18335 and b[50] n2685 ; n18591
g18336 and b[51] n2534 ; n18592
g18337 and n18591_not n18592_not ; n18593
g18338 and n18590_not n18593 ; n18594
g18339 and n2542_not n18594 ; n18595
g18340 and n9628_not n18594 ; n18596
g18341 and n18595_not n18596_not ; n18597
g18342 and a[26] n18597_not ; n18598
g18343 and a[26]_not n18597 ; n18599
g18344 and n18598_not n18599_not ; n18600
g18345 and n18589_not n18600_not ; n18601
g18346 and n18589 n18600 ; n18602
g18347 and n18601_not n18602_not ; n18603
g18348 and n18587_not n18603 ; n18604
g18349 and n18587_not n18604_not ; n18605
g18350 and n18603 n18604_not ; n18606
g18351 and n18605_not n18606_not ; n18607
g18352 and n18351_not n18607_not ; n18608
g18353 and n18351_not n18608_not ; n18609
g18354 and n18607_not n18608_not ; n18610
g18355 and n18609_not n18610_not ; n18611
g18356 and n18032_not n18293_not ; n18612
g18357 and b[58] n1627 ; n18613
g18358 and b[56] n1763 ; n18614
g18359 and b[57] n1622 ; n18615
g18360 and n18614_not n18615_not ; n18616
g18361 and n18613_not n18616 ; n18617
g18362 and n1630_not n18617 ; n18618
g18363 and n11436_not n18617 ; n18619
g18364 and n18618_not n18619_not ; n18620
g18365 and a[20] n18620_not ; n18621
g18366 and a[20]_not n18620 ; n18622
g18367 and n18621_not n18622_not ; n18623
g18368 and n18612_not n18623_not ; n18624
g18369 and n18612_not n18624_not ; n18625
g18370 and n18623_not n18624_not ; n18626
g18371 and n18625_not n18626_not ; n18627
g18372 and n18611_not n18627_not ; n18628
g18373 and n18611_not n18628_not ; n18629
g18374 and n18627_not n18628_not ; n18630
g18375 and n18629_not n18630_not ; n18631
g18376 and n18335_not n18631_not ; n18632
g18377 and n18335_not n18632_not ; n18633
g18378 and n18631_not n18632_not ; n18634
g18379 and n18633_not n18634_not ; n18635
g18380 and n17990_not n18001_not ; n18636
g18381 and n18301_not n18636_not ; n18637
g18382 and b[62] n1056 ; n18638
g18383 and b[63] n946 ; n18639
g18384 and n18638_not n18639_not ; n18640
g18385 and n954_not n18640 ; n18641
g18386 and n13800 n18640 ; n18642
g18387 and n18641_not n18642_not ; n18643
g18388 and a[14] n18643_not ; n18644
g18389 and a[14]_not n18643 ; n18645
g18390 and n18644_not n18645_not ; n18646
g18391 and n18637_not n18646_not ; n18647
g18392 and n18637_not n18647_not ; n18648
g18393 and n18646_not n18647_not ; n18649
g18394 and n18648_not n18649_not ; n18650
g18395 and n18635_not n18650_not ; n18651
g18396 and n18635 n18649_not ; n18652
g18397 and n18648_not n18652 ; n18653
g18398 and n18651_not n18653_not ; n18654
g18399 and n18319_not n18654 ; n18655
g18400 and n18319_not n18655_not ; n18656
g18401 and n18654 n18655_not ; n18657
g18402 and n18656_not n18657_not ; n18658
g18403 and n18317_not n18658_not ; n18659
g18404 and n18317 n18657_not ; n18660
g18405 and n18656_not n18660 ; n18661
g18406 and n18659_not n18661_not ; f[76]
g18407 and n18655_not n18659_not ; n18663
g18408 and n18647_not n18651_not ; n18664
g18409 and n18332_not n18632_not ; n18665
g18410 and b[63] n1056 ; n18666
g18411 and n954 n13797 ; n18667
g18412 and n18666_not n18667_not ; n18668
g18413 and a[14] n18668_not ; n18669
g18414 and a[14] n18669_not ; n18670
g18415 and n18668_not n18669_not ; n18671
g18416 and n18670_not n18671_not ; n18672
g18417 and n18665_not n18672_not ; n18673
g18418 and n18665_not n18673_not ; n18674
g18419 and n18672_not n18673_not ; n18675
g18420 and n18674_not n18675_not ; n18676
g18421 and b[59] n1627 ; n18677
g18422 and b[57] n1763 ; n18678
g18423 and b[58] n1622 ; n18679
g18424 and n18678_not n18679_not ; n18680
g18425 and n18677_not n18680 ; n18681
g18426 and n1630 n12179 ; n18682
g18427 and n18681 n18682_not ; n18683
g18428 and a[20] n18683_not ; n18684
g18429 and a[20] n18684_not ; n18685
g18430 and n18683_not n18684_not ; n18686
g18431 and n18685_not n18686_not ; n18687
g18432 and n18348_not n18608_not ; n18688
g18433 and n18687 n18688 ; n18689
g18434 and n18687_not n18688_not ; n18690
g18435 and n18689_not n18690_not ; n18691
g18436 and b[56] n2048 ; n18692
g18437 and b[54] n2198 ; n18693
g18438 and b[55] n2043 ; n18694
g18439 and n18693_not n18694_not ; n18695
g18440 and n18692_not n18695 ; n18696
g18441 and n2051 n10708 ; n18697
g18442 and n18696 n18697_not ; n18698
g18443 and a[23] n18698_not ; n18699
g18444 and a[23] n18699_not ; n18700
g18445 and n18698_not n18699_not ; n18701
g18446 and n18700_not n18701_not ; n18702
g18447 and n18601_not n18604_not ; n18703
g18448 and n18702 n18703 ; n18704
g18449 and n18702_not n18703_not ; n18705
g18450 and n18704_not n18705_not ; n18706
g18451 and b[53] n2539 ; n18707
g18452 and b[51] n2685 ; n18708
g18453 and b[52] n2534 ; n18709
g18454 and n18708_not n18709_not ; n18710
g18455 and n18707_not n18710 ; n18711
g18456 and n2542 n9972 ; n18712
g18457 and n18711 n18712_not ; n18713
g18458 and a[26] n18713_not ; n18714
g18459 and a[26] n18714_not ; n18715
g18460 and n18713_not n18714_not ; n18716
g18461 and n18715_not n18716_not ; n18717
g18462 and n18364_not n18584_not ; n18718
g18463 and n18717 n18718 ; n18719
g18464 and n18717_not n18718_not ; n18720
g18465 and n18719_not n18720_not ; n18721
g18466 and n18557_not n18560_not ; n18722
g18467 and b[47] n3638 ; n18723
g18468 and b[45] n3843 ; n18724
g18469 and b[46] n3633 ; n18725
g18470 and n18724_not n18725_not ; n18726
g18471 and n18723_not n18726 ; n18727
g18472 and n3641_not n18727 ; n18728
g18473 and n7703_not n18727 ; n18729
g18474 and n18728_not n18729_not ; n18730
g18475 and a[32] n18730_not ; n18731
g18476 and a[32]_not n18730 ; n18732
g18477 and n18731_not n18732_not ; n18733
g18478 and n18722_not n18733_not ; n18734
g18479 and n18722 n18733 ; n18735
g18480 and n18734_not n18735_not ; n18736
g18481 and b[44] n4287 ; n18737
g18482 and b[42] n4532 ; n18738
g18483 and b[43] n4282 ; n18739
g18484 and n18738_not n18739_not ; n18740
g18485 and n18737_not n18740 ; n18741
g18486 and n4290 n7072 ; n18742
g18487 and n18741 n18742_not ; n18743
g18488 and a[35] n18743_not ; n18744
g18489 and a[35] n18744_not ; n18745
g18490 and n18743_not n18744_not ; n18746
g18491 and n18745_not n18746_not ; n18747
g18492 and n18549_not n18553_not ; n18748
g18493 and b[41] n5035 ; n18749
g18494 and b[39] n5277 ; n18750
g18495 and b[40] n5030 ; n18751
g18496 and n18750_not n18751_not ; n18752
g18497 and n18749_not n18752 ; n18753
g18498 and n5038 n6219 ; n18754
g18499 and n18753 n18754_not ; n18755
g18500 and a[38] n18755_not ; n18756
g18501 and a[38] n18756_not ; n18757
g18502 and n18755_not n18756_not ; n18758
g18503 and n18757_not n18758_not ; n18759
g18504 and n18541_not n18545_not ; n18760
g18505 and n18527_not n18531_not ; n18761
g18506 and n18492_not n18505_not ; n18762
g18507 and b[26] n9339 ; n18763
g18508 and b[24] n9732 ; n18764
g18509 and b[25] n9334 ; n18765
g18510 and n18764_not n18765_not ; n18766
g18511 and n18763_not n18766 ; n18767
g18512 and n2813 n9342 ; n18768
g18513 and n18767 n18768_not ; n18769
g18514 and a[53] n18769_not ; n18770
g18515 and a[53] n18770_not ; n18771
g18516 and n18769_not n18770_not ; n18772
g18517 and n18771_not n18772_not ; n18773
g18518 and n18473_not n18486_not ; n18774
g18519 and n18437_not n18448_not ; n18775
g18520 and n18434_not n18775_not ; n18776
g18521 and b[13] n13903 ; n18777
g18522 and b[14] n13488_not ; n18778
g18523 and n18777_not n18778_not ; n18779
g18524 and n18431 n18779_not ; n18780
g18525 and n18431_not n18779 ; n18781
g18526 and n18780_not n18781_not ; n18782
g18527 and b[17] n12668 ; n18783
g18528 and b[15] n13047 ; n18784
g18529 and b[16] n12663 ; n18785
g18530 and n18784_not n18785_not ; n18786
g18531 and n18783_not n18786 ; n18787
g18532 and n12671_not n18787 ; n18788
g18533 and n1356_not n18787 ; n18789
g18534 and n18788_not n18789_not ; n18790
g18535 and a[62] n18790_not ; n18791
g18536 and a[62]_not n18790 ; n18792
g18537 and n18791_not n18792_not ; n18793
g18538 and n18782 n18793_not ; n18794
g18539 and n18782_not n18793 ; n18795
g18540 and n18794_not n18795_not ; n18796
g18541 and n18776_not n18796 ; n18797
g18542 and n18776 n18796_not ; n18798
g18543 and n18797_not n18798_not ; n18799
g18544 and b[20] n11531 ; n18800
g18545 and b[18] n11896 ; n18801
g18546 and b[19] n11526 ; n18802
g18547 and n18801_not n18802_not ; n18803
g18548 and n18800_not n18803 ; n18804
g18549 and n1846 n11534 ; n18805
g18550 and n18804 n18805_not ; n18806
g18551 and a[59] n18806_not ; n18807
g18552 and a[59] n18807_not ; n18808
g18553 and n18806_not n18807_not ; n18809
g18554 and n18808_not n18809_not ; n18810
g18555 and n18799 n18810_not ; n18811
g18556 and n18799 n18811_not ; n18812
g18557 and n18810_not n18811_not ; n18813
g18558 and n18812_not n18813_not ; n18814
g18559 and n18454_not n18467_not ; n18815
g18560 and n18814 n18815 ; n18816
g18561 and n18814_not n18815_not ; n18817
g18562 and n18816_not n18817_not ; n18818
g18563 and b[23] n10426 ; n18819
g18564 and b[21] n10796 ; n18820
g18565 and b[22] n10421 ; n18821
g18566 and n18820_not n18821_not ; n18822
g18567 and n18819_not n18822 ; n18823
g18568 and n2300 n10429 ; n18824
g18569 and n18823 n18824_not ; n18825
g18570 and a[56] n18825_not ; n18826
g18571 and a[56] n18826_not ; n18827
g18572 and n18825_not n18826_not ; n18828
g18573 and n18827_not n18828_not ; n18829
g18574 and n18818_not n18829 ; n18830
g18575 and n18818 n18829_not ; n18831
g18576 and n18830_not n18831_not ; n18832
g18577 and n18774_not n18832 ; n18833
g18578 and n18774 n18832_not ; n18834
g18579 and n18833_not n18834_not ; n18835
g18580 and n18773_not n18835 ; n18836
g18581 and n18773 n18835_not ; n18837
g18582 and n18836_not n18837_not ; n18838
g18583 and n18762_not n18838 ; n18839
g18584 and n18762 n18838_not ; n18840
g18585 and n18839_not n18840_not ; n18841
g18586 and b[29] n8362 ; n18842
g18587 and b[27] n8715 ; n18843
g18588 and b[28] n8357 ; n18844
g18589 and n18843_not n18844_not ; n18845
g18590 and n18842_not n18845 ; n18846
g18591 and n3383 n8365 ; n18847
g18592 and n18846 n18847_not ; n18848
g18593 and a[50] n18848_not ; n18849
g18594 and a[50] n18849_not ; n18850
g18595 and n18848_not n18849_not ; n18851
g18596 and n18850_not n18851_not ; n18852
g18597 and n18841 n18852_not ; n18853
g18598 and n18841 n18853_not ; n18854
g18599 and n18852_not n18853_not ; n18855
g18600 and n18854_not n18855_not ; n18856
g18601 and n18511_not n18525_not ; n18857
g18602 and n18856_not n18857_not ; n18858
g18603 and n18856_not n18858_not ; n18859
g18604 and n18857_not n18858_not ; n18860
g18605 and n18859_not n18860_not ; n18861
g18606 and b[32] n7446 ; n18862
g18607 and b[30] n7787 ; n18863
g18608 and b[31] n7441 ; n18864
g18609 and n18863_not n18864_not ; n18865
g18610 and n18862_not n18865 ; n18866
g18611 and n4013 n7449 ; n18867
g18612 and n18866 n18867_not ; n18868
g18613 and a[47] n18868_not ; n18869
g18614 and a[47] n18869_not ; n18870
g18615 and n18868_not n18869_not ; n18871
g18616 and n18870_not n18871_not ; n18872
g18617 and n18861_not n18872 ; n18873
g18618 and n18861 n18872_not ; n18874
g18619 and n18873_not n18874_not ; n18875
g18620 and n18761 n18875 ; n18876
g18621 and n18761_not n18875_not ; n18877
g18622 and n18876_not n18877_not ; n18878
g18623 and b[35] n6595 ; n18879
g18624 and b[33] n6902 ; n18880
g18625 and b[34] n6590 ; n18881
g18626 and n18880_not n18881_not ; n18882
g18627 and n18879_not n18882 ; n18883
g18628 and n4696 n6598 ; n18884
g18629 and n18883 n18884_not ; n18885
g18630 and a[44] n18885_not ; n18886
g18631 and a[44] n18886_not ; n18887
g18632 and n18885_not n18886_not ; n18888
g18633 and n18887_not n18888_not ; n18889
g18634 and n18878 n18889_not ; n18890
g18635 and n18878 n18890_not ; n18891
g18636 and n18889_not n18890_not ; n18892
g18637 and n18891_not n18892_not ; n18893
g18638 and n18535_not n18538_not ; n18894
g18639 and n18893 n18894 ; n18895
g18640 and n18893_not n18894_not ; n18896
g18641 and n18895_not n18896_not ; n18897
g18642 and b[38] n5777 ; n18898
g18643 and b[36] n6059 ; n18899
g18644 and b[37] n5772 ; n18900
g18645 and n18899_not n18900_not ; n18901
g18646 and n18898_not n18901 ; n18902
g18647 and n5205 n5780 ; n18903
g18648 and n18902 n18903_not ; n18904
g18649 and a[41] n18904_not ; n18905
g18650 and a[41] n18905_not ; n18906
g18651 and n18904_not n18905_not ; n18907
g18652 and n18906_not n18907_not ; n18908
g18653 and n18897_not n18908 ; n18909
g18654 and n18897 n18908_not ; n18910
g18655 and n18909_not n18910_not ; n18911
g18656 and n18760_not n18911 ; n18912
g18657 and n18760 n18911_not ; n18913
g18658 and n18912_not n18913_not ; n18914
g18659 and n18759_not n18914 ; n18915
g18660 and n18759 n18914_not ; n18916
g18661 and n18915_not n18916_not ; n18917
g18662 and n18748_not n18917 ; n18918
g18663 and n18748 n18917_not ; n18919
g18664 and n18918_not n18919_not ; n18920
g18665 and n18747_not n18920 ; n18921
g18666 and n18747_not n18921_not ; n18922
g18667 and n18920 n18921_not ; n18923
g18668 and n18922_not n18923_not ; n18924
g18669 and n18736 n18924_not ; n18925
g18670 and n18736 n18925_not ; n18926
g18671 and n18924_not n18925_not ; n18927
g18672 and n18926_not n18927_not ; n18928
g18673 and n18576_not n18580_not ; n18929
g18674 and b[50] n3050 ; n18930
g18675 and b[48] n3243 ; n18931
g18676 and b[49] n3045 ; n18932
g18677 and n18931_not n18932_not ; n18933
g18678 and n18930_not n18933 ; n18934
g18679 and n3053_not n18934 ; n18935
g18680 and n8949_not n18934 ; n18936
g18681 and n18935_not n18936_not ; n18937
g18682 and a[29] n18937_not ; n18938
g18683 and a[29]_not n18937 ; n18939
g18684 and n18938_not n18939_not ; n18940
g18685 and n18929_not n18940_not ; n18941
g18686 and n18929 n18940 ; n18942
g18687 and n18941_not n18942_not ; n18943
g18688 and n18928_not n18943 ; n18944
g18689 and n18928_not n18944_not ; n18945
g18690 and n18943 n18944_not ; n18946
g18691 and n18945_not n18946_not ; n18947
g18692 and n18721 n18947_not ; n18948
g18693 and n18721 n18948_not ; n18949
g18694 and n18947_not n18948_not ; n18950
g18695 and n18949_not n18950_not ; n18951
g18696 and n18706 n18951_not ; n18952
g18697 and n18706_not n18951 ; n18953
g18698 and n18691 n18953_not ; n18954
g18699 and n18952_not n18954 ; n18955
g18700 and n18691 n18955_not ; n18956
g18701 and n18953_not n18955_not ; n18957
g18702 and n18952_not n18957 ; n18958
g18703 and n18956_not n18958_not ; n18959
g18704 and n18624_not n18628_not ; n18960
g18705 and b[62] n1302 ; n18961
g18706 and b[60] n1391 ; n18962
g18707 and b[61] n1297 ; n18963
g18708 and n18962_not n18963_not ; n18964
g18709 and n18961_not n18964 ; n18965
g18710 and n1305_not n18965 ; n18966
g18711 and n13370_not n18965 ; n18967
g18712 and n18966_not n18967_not ; n18968
g18713 and a[17] n18968_not ; n18969
g18714 and a[17]_not n18968 ; n18970
g18715 and n18969_not n18970_not ; n18971
g18716 and n18960_not n18971_not ; n18972
g18717 and n18960_not n18972_not ; n18973
g18718 and n18971_not n18972_not ; n18974
g18719 and n18973_not n18974_not ; n18975
g18720 and n18959_not n18975_not ; n18976
g18721 and n18959 n18974_not ; n18977
g18722 and n18973_not n18977 ; n18978
g18723 and n18976_not n18978_not ; n18979
g18724 and n18676_not n18979 ; n18980
g18725 and n18676 n18979_not ; n18981
g18726 and n18980_not n18981_not ; n18982
g18727 and n18664_not n18982 ; n18983
g18728 and n18664 n18982_not ; n18984
g18729 and n18983_not n18984_not ; n18985
g18730 and n18663_not n18985 ; n18986
g18731 and n18663 n18985_not ; n18987
g18732 and n18986_not n18987_not ; f[77]
g18733 and n18972_not n18976_not ; n18989
g18734 and b[63] n1302 ; n18990
g18735 and b[61] n1391 ; n18991
g18736 and b[62] n1297 ; n18992
g18737 and n18991_not n18992_not ; n18993
g18738 and n18990_not n18993 ; n18994
g18739 and n1305 n13771 ; n18995
g18740 and n18994 n18995_not ; n18996
g18741 and a[17] n18996_not ; n18997
g18742 and a[17] n18997_not ; n18998
g18743 and n18996_not n18997_not ; n18999
g18744 and n18998_not n18999_not ; n19000
g18745 and n18989_not n19000_not ; n19001
g18746 and n18989_not n19001_not ; n19002
g18747 and n19000_not n19001_not ; n19003
g18748 and n19002_not n19003_not ; n19004
g18749 and b[60] n1627 ; n19005
g18750 and b[58] n1763 ; n19006
g18751 and b[59] n1622 ; n19007
g18752 and n19006_not n19007_not ; n19008
g18753 and n19005_not n19008 ; n19009
g18754 and n1630 n12211 ; n19010
g18755 and n19009 n19010_not ; n19011
g18756 and a[20] n19011_not ; n19012
g18757 and a[20] n19012_not ; n19013
g18758 and n19011_not n19012_not ; n19014
g18759 and n19013_not n19014_not ; n19015
g18760 and n18690_not n18955_not ; n19016
g18761 and n19015 n19016 ; n19017
g18762 and n19015_not n19016_not ; n19018
g18763 and n19017_not n19018_not ; n19019
g18764 and n18705_not n18952_not ; n19020
g18765 and b[57] n2048 ; n19021
g18766 and b[55] n2198 ; n19022
g18767 and b[56] n2043 ; n19023
g18768 and n19022_not n19023_not ; n19024
g18769 and n19021_not n19024 ; n19025
g18770 and n2051 n11410 ; n19026
g18771 and n19025 n19026_not ; n19027
g18772 and a[23] n19027_not ; n19028
g18773 and a[23] n19028_not ; n19029
g18774 and n19027_not n19028_not ; n19030
g18775 and n19029_not n19030_not ; n19031
g18776 and n19020_not n19031 ; n19032
g18777 and n19020 n19031_not ; n19033
g18778 and n19032_not n19033_not ; n19034
g18779 and b[54] n2539 ; n19035
g18780 and b[52] n2685 ; n19036
g18781 and b[53] n2534 ; n19037
g18782 and n19036_not n19037_not ; n19038
g18783 and n19035_not n19038 ; n19039
g18784 and n2542 n9998 ; n19040
g18785 and n19039 n19040_not ; n19041
g18786 and a[26] n19041_not ; n19042
g18787 and a[26] n19042_not ; n19043
g18788 and n19041_not n19042_not ; n19044
g18789 and n19043_not n19044_not ; n19045
g18790 and n18720_not n18948_not ; n19046
g18791 and n19045 n19046 ; n19047
g18792 and n19045_not n19046_not ; n19048
g18793 and n19047_not n19048_not ; n19049
g18794 and b[51] n3050 ; n19050
g18795 and b[49] n3243 ; n19051
g18796 and b[50] n3045 ; n19052
g18797 and n19051_not n19052_not ; n19053
g18798 and n19050_not n19053 ; n19054
g18799 and n3053 n8976 ; n19055
g18800 and n19054 n19055_not ; n19056
g18801 and a[29] n19056_not ; n19057
g18802 and a[29] n19057_not ; n19058
g18803 and n19056_not n19057_not ; n19059
g18804 and n19058_not n19059_not ; n19060
g18805 and n18941_not n18944_not ; n19061
g18806 and n19060 n19061 ; n19062
g18807 and n19060_not n19061_not ; n19063
g18808 and n19062_not n19063_not ; n19064
g18809 and n18912_not n18915_not ; n19065
g18810 and n18896_not n18910_not ; n19066
g18811 and n18877_not n18890_not ; n19067
g18812 and n18861_not n18872_not ; n19068
g18813 and n18858_not n19068_not ; n19069
g18814 and n18817_not n18831_not ; n19070
g18815 and b[14] n13903 ; n19071
g18816 and b[15] n13488_not ; n19072
g18817 and n19071_not n19072_not ; n19073
g18818 and a[14]_not n19073_not ; n19074
g18819 and a[14]_not n19074_not ; n19075
g18820 and n19073_not n19074_not ; n19076
g18821 and n19075_not n19076_not ; n19077
g18822 and n18431_not n19077_not ; n19078
g18823 and n18431_not n19078_not ; n19079
g18824 and n19077_not n19078_not ; n19080
g18825 and n19079_not n19080_not ; n19081
g18826 and b[18] n12668 ; n19082
g18827 and b[16] n13047 ; n19083
g18828 and b[17] n12663 ; n19084
g18829 and n19083_not n19084_not ; n19085
g18830 and n19082_not n19085 ; n19086
g18831 and n1566 n12671 ; n19087
g18832 and n19086 n19087_not ; n19088
g18833 and a[62] n19088_not ; n19089
g18834 and a[62] n19089_not ; n19090
g18835 and n19088_not n19089_not ; n19091
g18836 and n19090_not n19091_not ; n19092
g18837 and n19081_not n19092_not ; n19093
g18838 and n19081_not n19093_not ; n19094
g18839 and n19092_not n19093_not ; n19095
g18840 and n19094_not n19095_not ; n19096
g18841 and n18780_not n18794_not ; n19097
g18842 and n19096 n19097 ; n19098
g18843 and n19096_not n19097_not ; n19099
g18844 and n19098_not n19099_not ; n19100
g18845 and b[21] n11531 ; n19101
g18846 and b[19] n11896 ; n19102
g18847 and b[20] n11526 ; n19103
g18848 and n19102_not n19103_not ; n19104
g18849 and n19101_not n19104 ; n19105
g18850 and n1984 n11534 ; n19106
g18851 and n19105 n19106_not ; n19107
g18852 and a[59] n19107_not ; n19108
g18853 and a[59] n19108_not ; n19109
g18854 and n19107_not n19108_not ; n19110
g18855 and n19109_not n19110_not ; n19111
g18856 and n19100 n19111_not ; n19112
g18857 and n19100 n19112_not ; n19113
g18858 and n19111_not n19112_not ; n19114
g18859 and n19113_not n19114_not ; n19115
g18860 and n18797_not n18811_not ; n19116
g18861 and n19115 n19116 ; n19117
g18862 and n19115_not n19116_not ; n19118
g18863 and n19117_not n19118_not ; n19119
g18864 and b[24] n10426 ; n19120
g18865 and b[22] n10796 ; n19121
g18866 and b[23] n10421 ; n19122
g18867 and n19121_not n19122_not ; n19123
g18868 and n19120_not n19123 ; n19124
g18869 and n2458 n10429 ; n19125
g18870 and n19124 n19125_not ; n19126
g18871 and a[56] n19126_not ; n19127
g18872 and a[56] n19127_not ; n19128
g18873 and n19126_not n19127_not ; n19129
g18874 and n19128_not n19129_not ; n19130
g18875 and n19119 n19130_not ; n19131
g18876 and n19119_not n19130 ; n19132
g18877 and n19070_not n19132_not ; n19133
g18878 and n19131_not n19133 ; n19134
g18879 and n19070_not n19134_not ; n19135
g18880 and n19131_not n19134_not ; n19136
g18881 and n19132_not n19136 ; n19137
g18882 and n19135_not n19137_not ; n19138
g18883 and b[27] n9339 ; n19139
g18884 and b[25] n9732 ; n19140
g18885 and b[26] n9334 ; n19141
g18886 and n19140_not n19141_not ; n19142
g18887 and n19139_not n19142 ; n19143
g18888 and n2990 n9342 ; n19144
g18889 and n19143 n19144_not ; n19145
g18890 and a[53] n19145_not ; n19146
g18891 and a[53] n19146_not ; n19147
g18892 and n19145_not n19146_not ; n19148
g18893 and n19147_not n19148_not ; n19149
g18894 and n19138_not n19149_not ; n19150
g18895 and n19138_not n19150_not ; n19151
g18896 and n19149_not n19150_not ; n19152
g18897 and n19151_not n19152_not ; n19153
g18898 and n18833_not n18836_not ; n19154
g18899 and n19153 n19154 ; n19155
g18900 and n19153_not n19154_not ; n19156
g18901 and n19155_not n19156_not ; n19157
g18902 and b[30] n8362 ; n19158
g18903 and b[28] n8715 ; n19159
g18904 and b[29] n8357 ; n19160
g18905 and n19159_not n19160_not ; n19161
g18906 and n19158_not n19161 ; n19162
g18907 and n3577 n8365 ; n19163
g18908 and n19162 n19163_not ; n19164
g18909 and a[50] n19164_not ; n19165
g18910 and a[50] n19165_not ; n19166
g18911 and n19164_not n19165_not ; n19167
g18912 and n19166_not n19167_not ; n19168
g18913 and n19157 n19168_not ; n19169
g18914 and n19157 n19169_not ; n19170
g18915 and n19168_not n19169_not ; n19171
g18916 and n19170_not n19171_not ; n19172
g18917 and n18839_not n18853_not ; n19173
g18918 and n19172 n19173 ; n19174
g18919 and n19172_not n19173_not ; n19175
g18920 and n19174_not n19175_not ; n19176
g18921 and b[33] n7446 ; n19177
g18922 and b[31] n7787 ; n19178
g18923 and b[32] n7441 ; n19179
g18924 and n19178_not n19179_not ; n19180
g18925 and n19177_not n19180 ; n19181
g18926 and n4223 n7449 ; n19182
g18927 and n19181 n19182_not ; n19183
g18928 and a[47] n19183_not ; n19184
g18929 and a[47] n19184_not ; n19185
g18930 and n19183_not n19184_not ; n19186
g18931 and n19185_not n19186_not ; n19187
g18932 and n19176 n19187_not ; n19188
g18933 and n19176 n19188_not ; n19189
g18934 and n19187_not n19188_not ; n19190
g18935 and n19189_not n19190_not ; n19191
g18936 and n19069_not n19191 ; n19192
g18937 and n19069 n19191_not ; n19193
g18938 and n19192_not n19193_not ; n19194
g18939 and b[36] n6595 ; n19195
g18940 and b[34] n6902 ; n19196
g18941 and b[35] n6590 ; n19197
g18942 and n19196_not n19197_not ; n19198
g18943 and n19195_not n19198 ; n19199
g18944 and n4922 n6598 ; n19200
g18945 and n19199 n19200_not ; n19201
g18946 and a[44] n19201_not ; n19202
g18947 and a[44] n19202_not ; n19203
g18948 and n19201_not n19202_not ; n19204
g18949 and n19203_not n19204_not ; n19205
g18950 and n19194_not n19205_not ; n19206
g18951 and n19194 n19205 ; n19207
g18952 and n19206_not n19207_not ; n19208
g18953 and n19067 n19208_not ; n19209
g18954 and n19067_not n19208 ; n19210
g18955 and n19209_not n19210_not ; n19211
g18956 and b[39] n5777 ; n19212
g18957 and b[37] n6059 ; n19213
g18958 and b[38] n5772 ; n19214
g18959 and n19213_not n19214_not ; n19215
g18960 and n19212_not n19215 ; n19216
g18961 and n5451 n5780 ; n19217
g18962 and n19216 n19217_not ; n19218
g18963 and a[41] n19218_not ; n19219
g18964 and a[41] n19219_not ; n19220
g18965 and n19218_not n19219_not ; n19221
g18966 and n19220_not n19221_not ; n19222
g18967 and n19211 n19222_not ; n19223
g18968 and n19211 n19223_not ; n19224
g18969 and n19222_not n19223_not ; n19225
g18970 and n19224_not n19225_not ; n19226
g18971 and n19066_not n19226 ; n19227
g18972 and n19066 n19226_not ; n19228
g18973 and n19227_not n19228_not ; n19229
g18974 and b[42] n5035 ; n19230
g18975 and b[40] n5277 ; n19231
g18976 and b[41] n5030 ; n19232
g18977 and n19231_not n19232_not ; n19233
g18978 and n19230_not n19233 ; n19234
g18979 and n5038 n6489 ; n19235
g18980 and n19234 n19235_not ; n19236
g18981 and a[38] n19236_not ; n19237
g18982 and a[38] n19237_not ; n19238
g18983 and n19236_not n19237_not ; n19239
g18984 and n19238_not n19239_not ; n19240
g18985 and n19229_not n19240_not ; n19241
g18986 and n19229 n19240 ; n19242
g18987 and n19241_not n19242_not ; n19243
g18988 and n19065 n19243_not ; n19244
g18989 and n19065_not n19243 ; n19245
g18990 and n19244_not n19245_not ; n19246
g18991 and b[45] n4287 ; n19247
g18992 and b[43] n4532 ; n19248
g18993 and b[44] n4282 ; n19249
g18994 and n19248_not n19249_not ; n19250
g18995 and n19247_not n19250 ; n19251
g18996 and n4290 n7361 ; n19252
g18997 and n19251 n19252_not ; n19253
g18998 and a[35] n19253_not ; n19254
g18999 and a[35] n19254_not ; n19255
g19000 and n19253_not n19254_not ; n19256
g19001 and n19255_not n19256_not ; n19257
g19002 and n19246 n19257_not ; n19258
g19003 and n19246 n19258_not ; n19259
g19004 and n19257_not n19258_not ; n19260
g19005 and n19259_not n19260_not ; n19261
g19006 and n18918_not n18921_not ; n19262
g19007 and n19261 n19262 ; n19263
g19008 and n19261_not n19262_not ; n19264
g19009 and n19263_not n19264_not ; n19265
g19010 and n18734_not n18925_not ; n19266
g19011 and b[48] n3638 ; n19267
g19012 and b[46] n3843 ; n19268
g19013 and b[47] n3633 ; n19269
g19014 and n19268_not n19269_not ; n19270
g19015 and n19267_not n19270 ; n19271
g19016 and n3641 n8009 ; n19272
g19017 and n19271 n19272_not ; n19273
g19018 and a[32] n19273_not ; n19274
g19019 and a[32] n19274_not ; n19275
g19020 and n19273_not n19274_not ; n19276
g19021 and n19275_not n19276_not ; n19277
g19022 and n19266_not n19277_not ; n19278
g19023 and n19266_not n19278_not ; n19279
g19024 and n19277_not n19278_not ; n19280
g19025 and n19279_not n19280_not ; n19281
g19026 and n19265 n19281_not ; n19282
g19027 and n19265_not n19281 ; n19283
g19028 and n19064 n19283_not ; n19284
g19029 and n19282_not n19284 ; n19285
g19030 and n19064 n19285_not ; n19286
g19031 and n19283_not n19285_not ; n19287
g19032 and n19282_not n19287 ; n19288
g19033 and n19286_not n19288_not ; n19289
g19034 and n19049 n19289_not ; n19290
g19035 and n19049_not n19289 ; n19291
g19036 and n19034_not n19291_not ; n19292
g19037 and n19290_not n19292 ; n19293
g19038 and n19034_not n19293_not ; n19294
g19039 and n19291_not n19293_not ; n19295
g19040 and n19290_not n19295 ; n19296
g19041 and n19294_not n19296_not ; n19297
g19042 and n19019 n19297_not ; n19298
g19043 and n19019_not n19297 ; n19299
g19044 and n19004_not n19299_not ; n19300
g19045 and n19298_not n19300 ; n19301
g19046 and n19004_not n19301_not ; n19302
g19047 and n19299_not n19301_not ; n19303
g19048 and n19298_not n19303 ; n19304
g19049 and n19302_not n19304_not ; n19305
g19050 and n18673_not n18980_not ; n19306
g19051 and n19305 n19306 ; n19307
g19052 and n19305_not n19306_not ; n19308
g19053 and n19307_not n19308_not ; n19309
g19054 and n18983_not n18986_not ; n19310
g19055 and n19309 n19310_not ; n19311
g19056 and n19309_not n19310 ; n19312
g19057 and n19311_not n19312_not ; f[78]
g19058 and n19018_not n19298_not ; n19314
g19059 and b[62] n1391 ; n19315
g19060 and b[63] n1297 ; n19316
g19061 and n19315_not n19316_not ; n19317
g19062 and n1305_not n19317 ; n19318
g19063 and n13800 n19317 ; n19319
g19064 and n19318_not n19319_not ; n19320
g19065 and a[17] n19320_not ; n19321
g19066 and a[17]_not n19320 ; n19322
g19067 and n19321_not n19322_not ; n19323
g19068 and n19314_not n19323_not ; n19324
g19069 and n19314 n19323 ; n19325
g19070 and n19324_not n19325_not ; n19326
g19071 and b[61] n1627 ; n19327
g19072 and b[59] n1763 ; n19328
g19073 and b[60] n1622 ; n19329
g19074 and n19328_not n19329_not ; n19330
g19075 and n19327_not n19330 ; n19331
g19076 and n1630 n12969 ; n19332
g19077 and n19331 n19332_not ; n19333
g19078 and a[20] n19333_not ; n19334
g19079 and a[20] n19334_not ; n19335
g19080 and n19333_not n19334_not ; n19336
g19081 and n19335_not n19336_not ; n19337
g19082 and n19020_not n19031_not ; n19338
g19083 and n19293_not n19338_not ; n19339
g19084 and n19337 n19339 ; n19340
g19085 and n19337_not n19339_not ; n19341
g19086 and n19340_not n19341_not ; n19342
g19087 and n19048_not n19290_not ; n19343
g19088 and b[58] n2048 ; n19344
g19089 and b[56] n2198 ; n19345
g19090 and b[57] n2043 ; n19346
g19091 and n19345_not n19346_not ; n19347
g19092 and n19344_not n19347 ; n19348
g19093 and n2051_not n19348 ; n19349
g19094 and n11436_not n19348 ; n19350
g19095 and n19349_not n19350_not ; n19351
g19096 and a[23] n19351_not ; n19352
g19097 and a[23]_not n19351 ; n19353
g19098 and n19352_not n19353_not ; n19354
g19099 and n19343_not n19354_not ; n19355
g19100 and n19343 n19354 ; n19356
g19101 and n19355_not n19356_not ; n19357
g19102 and b[55] n2539 ; n19358
g19103 and b[53] n2685 ; n19359
g19104 and b[54] n2534 ; n19360
g19105 and n19359_not n19360_not ; n19361
g19106 and n19358_not n19361 ; n19362
g19107 and n2542 n10684 ; n19363
g19108 and n19362 n19363_not ; n19364
g19109 and a[26] n19364_not ; n19365
g19110 and a[26] n19365_not ; n19366
g19111 and n19364_not n19365_not ; n19367
g19112 and n19366_not n19367_not ; n19368
g19113 and n19063_not n19285_not ; n19369
g19114 and n19368 n19369 ; n19370
g19115 and n19368_not n19369_not ; n19371
g19116 and n19370_not n19371_not ; n19372
g19117 and b[52] n3050 ; n19373
g19118 and b[50] n3243 ; n19374
g19119 and b[51] n3045 ; n19375
g19120 and n19374_not n19375_not ; n19376
g19121 and n19373_not n19376 ; n19377
g19122 and n3053 n9628 ; n19378
g19123 and n19377 n19378_not ; n19379
g19124 and a[29] n19379_not ; n19380
g19125 and a[29] n19380_not ; n19381
g19126 and n19379_not n19380_not ; n19382
g19127 and n19381_not n19382_not ; n19383
g19128 and n19278_not n19282_not ; n19384
g19129 and n19383_not n19384_not ; n19385
g19130 and n19383_not n19385_not ; n19386
g19131 and n19384_not n19385_not ; n19387
g19132 and n19386_not n19387_not ; n19388
g19133 and b[49] n3638 ; n19389
g19134 and b[47] n3843 ; n19390
g19135 and b[48] n3633 ; n19391
g19136 and n19390_not n19391_not ; n19392
g19137 and n19389_not n19392 ; n19393
g19138 and n3641 n8625 ; n19394
g19139 and n19393 n19394_not ; n19395
g19140 and a[32] n19395_not ; n19396
g19141 and a[32] n19396_not ; n19397
g19142 and n19395_not n19396_not ; n19398
g19143 and n19397_not n19398_not ; n19399
g19144 and n19258_not n19264_not ; n19400
g19145 and n19399 n19400 ; n19401
g19146 and n19399_not n19400_not ; n19402
g19147 and n19401_not n19402_not ; n19403
g19148 and b[43] n5035 ; n19404
g19149 and b[41] n5277 ; n19405
g19150 and b[42] n5030 ; n19406
g19151 and n19405_not n19406_not ; n19407
g19152 and n19404_not n19407 ; n19408
g19153 and n5038 n6515 ; n19409
g19154 and n19408 n19409_not ; n19410
g19155 and a[38] n19410_not ; n19411
g19156 and a[38] n19411_not ; n19412
g19157 and n19410_not n19411_not ; n19413
g19158 and n19412_not n19413_not ; n19414
g19159 and n19066_not n19226_not ; n19415
g19160 and n19223_not n19415_not ; n19416
g19161 and b[40] n5777 ; n19417
g19162 and b[38] n6059 ; n19418
g19163 and b[39] n5772 ; n19419
g19164 and n19418_not n19419_not ; n19420
g19165 and n19417_not n19420 ; n19421
g19166 and n5780 n5955 ; n19422
g19167 and n19421 n19422_not ; n19423
g19168 and a[41] n19423_not ; n19424
g19169 and a[41] n19424_not ; n19425
g19170 and n19423_not n19424_not ; n19426
g19171 and n19425_not n19426_not ; n19427
g19172 and n19206_not n19210_not ; n19428
g19173 and b[37] n6595 ; n19429
g19174 and b[35] n6902 ; n19430
g19175 and b[36] n6590 ; n19431
g19176 and n19430_not n19431_not ; n19432
g19177 and n19429_not n19432 ; n19433
g19178 and n5181 n6598 ; n19434
g19179 and n19433 n19434_not ; n19435
g19180 and a[44] n19435_not ; n19436
g19181 and a[44] n19436_not ; n19437
g19182 and n19435_not n19436_not ; n19438
g19183 and n19437_not n19438_not ; n19439
g19184 and n19069_not n19191_not ; n19440
g19185 and n19188_not n19440_not ; n19441
g19186 and b[31] n8362 ; n19442
g19187 and b[29] n8715 ; n19443
g19188 and b[30] n8357 ; n19444
g19189 and n19443_not n19444_not ; n19445
g19190 and n19442_not n19445 ; n19446
g19191 and n3796 n8365 ; n19447
g19192 and n19446 n19447_not ; n19448
g19193 and a[50] n19448_not ; n19449
g19194 and a[50] n19449_not ; n19450
g19195 and n19448_not n19449_not ; n19451
g19196 and n19450_not n19451_not ; n19452
g19197 and n19093_not n19099_not ; n19453
g19198 and b[15] n13903 ; n19454
g19199 and b[16] n13488_not ; n19455
g19200 and n19454_not n19455_not ; n19456
g19201 and n19074_not n19078_not ; n19457
g19202 and n19456_not n19457 ; n19458
g19203 and n19456 n19457_not ; n19459
g19204 and n19458_not n19459_not ; n19460
g19205 and b[19] n12668 ; n19461
g19206 and b[17] n13047 ; n19462
g19207 and b[18] n12663 ; n19463
g19208 and n19462_not n19463_not ; n19464
g19209 and n19461_not n19464 ; n19465
g19210 and n12671_not n19465 ; n19466
g19211 and n1708_not n19465 ; n19467
g19212 and n19466_not n19467_not ; n19468
g19213 and a[62] n19468_not ; n19469
g19214 and a[62]_not n19468 ; n19470
g19215 and n19469_not n19470_not ; n19471
g19216 and n19460 n19471_not ; n19472
g19217 and n19460_not n19471 ; n19473
g19218 and n19472_not n19473_not ; n19474
g19219 and n19453_not n19474 ; n19475
g19220 and n19453 n19474_not ; n19476
g19221 and n19475_not n19476_not ; n19477
g19222 and b[22] n11531 ; n19478
g19223 and b[20] n11896 ; n19479
g19224 and b[21] n11526 ; n19480
g19225 and n19479_not n19480_not ; n19481
g19226 and n19478_not n19481 ; n19482
g19227 and n2145 n11534 ; n19483
g19228 and n19482 n19483_not ; n19484
g19229 and a[59] n19484_not ; n19485
g19230 and a[59] n19485_not ; n19486
g19231 and n19484_not n19485_not ; n19487
g19232 and n19486_not n19487_not ; n19488
g19233 and n19477 n19488_not ; n19489
g19234 and n19477 n19489_not ; n19490
g19235 and n19488_not n19489_not ; n19491
g19236 and n19490_not n19491_not ; n19492
g19237 and n19112_not n19118_not ; n19493
g19238 and n19492 n19493 ; n19494
g19239 and n19492_not n19493_not ; n19495
g19240 and n19494_not n19495_not ; n19496
g19241 and b[25] n10426 ; n19497
g19242 and b[23] n10796 ; n19498
g19243 and b[24] n10421 ; n19499
g19244 and n19498_not n19499_not ; n19500
g19245 and n19497_not n19500 ; n19501
g19246 and n2485 n10429 ; n19502
g19247 and n19501 n19502_not ; n19503
g19248 and a[56] n19503_not ; n19504
g19249 and a[56] n19504_not ; n19505
g19250 and n19503_not n19504_not ; n19506
g19251 and n19505_not n19506_not ; n19507
g19252 and n19496 n19507_not ; n19508
g19253 and n19496 n19508_not ; n19509
g19254 and n19507_not n19508_not ; n19510
g19255 and n19509_not n19510_not ; n19511
g19256 and n19136_not n19511 ; n19512
g19257 and n19136 n19511_not ; n19513
g19258 and n19512_not n19513_not ; n19514
g19259 and b[28] n9339 ; n19515
g19260 and b[26] n9732 ; n19516
g19261 and b[27] n9334 ; n19517
g19262 and n19516_not n19517_not ; n19518
g19263 and n19515_not n19518 ; n19519
g19264 and n3189 n9342 ; n19520
g19265 and n19519 n19520_not ; n19521
g19266 and a[53] n19521_not ; n19522
g19267 and a[53] n19522_not ; n19523
g19268 and n19521_not n19522_not ; n19524
g19269 and n19523_not n19524_not ; n19525
g19270 and n19514 n19525 ; n19526
g19271 and n19514_not n19525_not ; n19527
g19272 and n19526_not n19527_not ; n19528
g19273 and n19150_not n19156_not ; n19529
g19274 and n19528 n19529_not ; n19530
g19275 and n19528_not n19529 ; n19531
g19276 and n19530_not n19531_not ; n19532
g19277 and n19452_not n19532 ; n19533
g19278 and n19532 n19533_not ; n19534
g19279 and n19452_not n19533_not ; n19535
g19280 and n19534_not n19535_not ; n19536
g19281 and n19169_not n19175_not ; n19537
g19282 and n19536 n19537 ; n19538
g19283 and n19536_not n19537_not ; n19539
g19284 and n19538_not n19539_not ; n19540
g19285 and b[34] n7446 ; n19541
g19286 and b[32] n7787 ; n19542
g19287 and b[33] n7441 ; n19543
g19288 and n19542_not n19543_not ; n19544
g19289 and n19541_not n19544 ; n19545
g19290 and n4466 n7449 ; n19546
g19291 and n19545 n19546_not ; n19547
g19292 and a[47] n19547_not ; n19548
g19293 and a[47] n19548_not ; n19549
g19294 and n19547_not n19548_not ; n19550
g19295 and n19549_not n19550_not ; n19551
g19296 and n19540_not n19551 ; n19552
g19297 and n19540 n19551_not ; n19553
g19298 and n19552_not n19553_not ; n19554
g19299 and n19441_not n19554 ; n19555
g19300 and n19441_not n19555_not ; n19556
g19301 and n19554 n19555_not ; n19557
g19302 and n19556_not n19557_not ; n19558
g19303 and n19439_not n19558_not ; n19559
g19304 and n19439 n19557_not ; n19560
g19305 and n19556_not n19560 ; n19561
g19306 and n19559_not n19561_not ; n19562
g19307 and n19428_not n19562 ; n19563
g19308 and n19428_not n19563_not ; n19564
g19309 and n19562 n19563_not ; n19565
g19310 and n19564_not n19565_not ; n19566
g19311 and n19427_not n19566_not ; n19567
g19312 and n19427 n19565_not ; n19568
g19313 and n19564_not n19568 ; n19569
g19314 and n19567_not n19569_not ; n19570
g19315 and n19416_not n19570 ; n19571
g19316 and n19416 n19570_not ; n19572
g19317 and n19571_not n19572_not ; n19573
g19318 and n19414_not n19573 ; n19574
g19319 and n19573 n19574_not ; n19575
g19320 and n19414_not n19574_not ; n19576
g19321 and n19575_not n19576_not ; n19577
g19322 and n19241_not n19245_not ; n19578
g19323 and n19577 n19578 ; n19579
g19324 and n19577_not n19578_not ; n19580
g19325 and n19579_not n19580_not ; n19581
g19326 and b[46] n4287 ; n19582
g19327 and b[44] n4532 ; n19583
g19328 and b[45] n4282 ; n19584
g19329 and n19583_not n19584_not ; n19585
g19330 and n19582_not n19585 ; n19586
g19331 and n4290 n7677 ; n19587
g19332 and n19586 n19587_not ; n19588
g19333 and a[35] n19588_not ; n19589
g19334 and a[35] n19589_not ; n19590
g19335 and n19588_not n19589_not ; n19591
g19336 and n19590_not n19591_not ; n19592
g19337 and n19581 n19592_not ; n19593
g19338 and n19581 n19593_not ; n19594
g19339 and n19592_not n19593_not ; n19595
g19340 and n19594_not n19595_not ; n19596
g19341 and n19403 n19596_not ; n19597
g19342 and n19403_not n19596 ; n19598
g19343 and n19388_not n19598_not ; n19599
g19344 and n19597_not n19599 ; n19600
g19345 and n19388_not n19600_not ; n19601
g19346 and n19598_not n19600_not ; n19602
g19347 and n19597_not n19602 ; n19603
g19348 and n19601_not n19603_not ; n19604
g19349 and n19372 n19604_not ; n19605
g19350 and n19372_not n19604 ; n19606
g19351 and n19357 n19606_not ; n19607
g19352 and n19605_not n19607 ; n19608
g19353 and n19357 n19608_not ; n19609
g19354 and n19606_not n19608_not ; n19610
g19355 and n19605_not n19610 ; n19611
g19356 and n19609_not n19611_not ; n19612
g19357 and n19342 n19612_not ; n19613
g19358 and n19342_not n19612 ; n19614
g19359 and n19326 n19614_not ; n19615
g19360 and n19613_not n19615 ; n19616
g19361 and n19326 n19616_not ; n19617
g19362 and n19614_not n19616_not ; n19618
g19363 and n19613_not n19618 ; n19619
g19364 and n19617_not n19619_not ; n19620
g19365 and n19001_not n19301_not ; n19621
g19366 and n19620 n19621 ; n19622
g19367 and n19620_not n19621_not ; n19623
g19368 and n19622_not n19623_not ; n19624
g19369 and n19308_not n19311_not ; n19625
g19370 and n19624 n19625_not ; n19626
g19371 and n19624_not n19625 ; n19627
g19372 and n19626_not n19627_not ; f[79]
g19373 and n19623_not n19626_not ; n19629
g19374 and n19324_not n19616_not ; n19630
g19375 and n19341_not n19613_not ; n19631
g19376 and b[63] n1391 ; n19632
g19377 and n1305 n13797 ; n19633
g19378 and n19632_not n19633_not ; n19634
g19379 and a[17] n19634_not ; n19635
g19380 and a[17] n19635_not ; n19636
g19381 and n19634_not n19635_not ; n19637
g19382 and n19636_not n19637_not ; n19638
g19383 and n19631_not n19638_not ; n19639
g19384 and n19631_not n19639_not ; n19640
g19385 and n19638_not n19639_not ; n19641
g19386 and n19640_not n19641_not ; n19642
g19387 and b[62] n1627 ; n19643
g19388 and b[60] n1763 ; n19644
g19389 and b[61] n1622 ; n19645
g19390 and n19644_not n19645_not ; n19646
g19391 and n19643_not n19646 ; n19647
g19392 and n1630 n13370 ; n19648
g19393 and n19647 n19648_not ; n19649
g19394 and a[20] n19649_not ; n19650
g19395 and a[20] n19650_not ; n19651
g19396 and n19649_not n19650_not ; n19652
g19397 and n19651_not n19652_not ; n19653
g19398 and n19355_not n19608_not ; n19654
g19399 and n19653 n19654 ; n19655
g19400 and n19653_not n19654_not ; n19656
g19401 and n19655_not n19656_not ; n19657
g19402 and b[59] n2048 ; n19658
g19403 and b[57] n2198 ; n19659
g19404 and b[58] n2043 ; n19660
g19405 and n19659_not n19660_not ; n19661
g19406 and n19658_not n19661 ; n19662
g19407 and n2051 n12179 ; n19663
g19408 and n19662 n19663_not ; n19664
g19409 and a[23] n19664_not ; n19665
g19410 and a[23] n19665_not ; n19666
g19411 and n19664_not n19665_not ; n19667
g19412 and n19666_not n19667_not ; n19668
g19413 and n19371_not n19605_not ; n19669
g19414 and n19668_not n19669_not ; n19670
g19415 and n19668_not n19670_not ; n19671
g19416 and n19669_not n19670_not ; n19672
g19417 and n19671_not n19672_not ; n19673
g19418 and b[56] n2539 ; n19674
g19419 and b[54] n2685 ; n19675
g19420 and b[55] n2534 ; n19676
g19421 and n19675_not n19676_not ; n19677
g19422 and n19674_not n19677 ; n19678
g19423 and n2542 n10708 ; n19679
g19424 and n19678 n19679_not ; n19680
g19425 and a[26] n19680_not ; n19681
g19426 and a[26] n19681_not ; n19682
g19427 and n19680_not n19681_not ; n19683
g19428 and n19682_not n19683_not ; n19684
g19429 and n19385_not n19600_not ; n19685
g19430 and n19684 n19685 ; n19686
g19431 and n19684_not n19685_not ; n19687
g19432 and n19686_not n19687_not ; n19688
g19433 and b[53] n3050 ; n19689
g19434 and b[51] n3243 ; n19690
g19435 and b[52] n3045 ; n19691
g19436 and n19690_not n19691_not ; n19692
g19437 and n19689_not n19692 ; n19693
g19438 and n3053 n9972 ; n19694
g19439 and n19693 n19694_not ; n19695
g19440 and a[29] n19695_not ; n19696
g19441 and a[29] n19696_not ; n19697
g19442 and n19695_not n19696_not ; n19698
g19443 and n19697_not n19698_not ; n19699
g19444 and n19402_not n19597_not ; n19700
g19445 and n19699_not n19700_not ; n19701
g19446 and n19699_not n19701_not ; n19702
g19447 and n19700_not n19701_not ; n19703
g19448 and n19702_not n19703_not ; n19704
g19449 and b[50] n3638 ; n19705
g19450 and b[48] n3843 ; n19706
g19451 and b[49] n3633 ; n19707
g19452 and n19706_not n19707_not ; n19708
g19453 and n19705_not n19708 ; n19709
g19454 and n3641 n8949 ; n19710
g19455 and n19709 n19710_not ; n19711
g19456 and a[32] n19711_not ; n19712
g19457 and a[32] n19712_not ; n19713
g19458 and n19711_not n19712_not ; n19714
g19459 and n19713_not n19714_not ; n19715
g19460 and n19580_not n19593_not ; n19716
g19461 and n19715 n19716 ; n19717
g19462 and n19715_not n19716_not ; n19718
g19463 and n19717_not n19718_not ; n19719
g19464 and n19571_not n19574_not ; n19720
g19465 and b[44] n5035 ; n19721
g19466 and b[42] n5277 ; n19722
g19467 and b[43] n5030 ; n19723
g19468 and n19722_not n19723_not ; n19724
g19469 and n19721_not n19724 ; n19725
g19470 and n5038 n7072 ; n19726
g19471 and n19725 n19726_not ; n19727
g19472 and a[38] n19727_not ; n19728
g19473 and a[38] n19728_not ; n19729
g19474 and n19727_not n19728_not ; n19730
g19475 and n19729_not n19730_not ; n19731
g19476 and n19563_not n19567_not ; n19732
g19477 and b[41] n5777 ; n19733
g19478 and b[39] n6059 ; n19734
g19479 and b[40] n5772 ; n19735
g19480 and n19734_not n19735_not ; n19736
g19481 and n19733_not n19736 ; n19737
g19482 and n5780 n6219 ; n19738
g19483 and n19737 n19738_not ; n19739
g19484 and a[41] n19739_not ; n19740
g19485 and a[41] n19740_not ; n19741
g19486 and n19739_not n19740_not ; n19742
g19487 and n19741_not n19742_not ; n19743
g19488 and n19555_not n19559_not ; n19744
g19489 and n19495_not n19508_not ; n19745
g19490 and b[26] n10426 ; n19746
g19491 and b[24] n10796 ; n19747
g19492 and b[25] n10421 ; n19748
g19493 and n19747_not n19748_not ; n19749
g19494 and n19746_not n19749 ; n19750
g19495 and n2813 n10429 ; n19751
g19496 and n19750 n19751_not ; n19752
g19497 and a[56] n19752_not ; n19753
g19498 and a[56] n19753_not ; n19754
g19499 and n19752_not n19753_not ; n19755
g19500 and n19754_not n19755_not ; n19756
g19501 and n19475_not n19489_not ; n19757
g19502 and b[20] n12668 ; n19758
g19503 and b[18] n13047 ; n19759
g19504 and b[19] n12663 ; n19760
g19505 and n19759_not n19760_not ; n19761
g19506 and n19758_not n19761 ; n19762
g19507 and n1846 n12671 ; n19763
g19508 and n19762 n19763_not ; n19764
g19509 and a[62] n19764_not ; n19765
g19510 and a[62] n19765_not ; n19766
g19511 and n19764_not n19765_not ; n19767
g19512 and n19766_not n19767_not ; n19768
g19513 and b[16] n13903 ; n19769
g19514 and b[17] n13488_not ; n19770
g19515 and n19769_not n19770_not ; n19771
g19516 and n19456 n19771_not ; n19772
g19517 and n19456_not n19771 ; n19773
g19518 and n19768_not n19773_not ; n19774
g19519 and n19772_not n19774 ; n19775
g19520 and n19768_not n19775_not ; n19776
g19521 and n19773_not n19775_not ; n19777
g19522 and n19772_not n19777 ; n19778
g19523 and n19776_not n19778_not ; n19779
g19524 and n19459_not n19472_not ; n19780
g19525 and n19779 n19780 ; n19781
g19526 and n19779_not n19780_not ; n19782
g19527 and n19781_not n19782_not ; n19783
g19528 and b[23] n11531 ; n19784
g19529 and b[21] n11896 ; n19785
g19530 and b[22] n11526 ; n19786
g19531 and n19785_not n19786_not ; n19787
g19532 and n19784_not n19787 ; n19788
g19533 and n2300 n11534 ; n19789
g19534 and n19788 n19789_not ; n19790
g19535 and a[59] n19790_not ; n19791
g19536 and a[59] n19791_not ; n19792
g19537 and n19790_not n19791_not ; n19793
g19538 and n19792_not n19793_not ; n19794
g19539 and n19783_not n19794 ; n19795
g19540 and n19783 n19794_not ; n19796
g19541 and n19795_not n19796_not ; n19797
g19542 and n19757_not n19797 ; n19798
g19543 and n19757 n19797_not ; n19799
g19544 and n19798_not n19799_not ; n19800
g19545 and n19756_not n19800 ; n19801
g19546 and n19756 n19800_not ; n19802
g19547 and n19801_not n19802_not ; n19803
g19548 and n19745_not n19803 ; n19804
g19549 and n19745 n19803_not ; n19805
g19550 and n19804_not n19805_not ; n19806
g19551 and b[29] n9339 ; n19807
g19552 and b[27] n9732 ; n19808
g19553 and b[28] n9334 ; n19809
g19554 and n19808_not n19809_not ; n19810
g19555 and n19807_not n19810 ; n19811
g19556 and n3383 n9342 ; n19812
g19557 and n19811 n19812_not ; n19813
g19558 and a[53] n19813_not ; n19814
g19559 and a[53] n19814_not ; n19815
g19560 and n19813_not n19814_not ; n19816
g19561 and n19815_not n19816_not ; n19817
g19562 and n19806 n19817_not ; n19818
g19563 and n19806 n19818_not ; n19819
g19564 and n19817_not n19818_not ; n19820
g19565 and n19819_not n19820_not ; n19821
g19566 and n19136_not n19511_not ; n19822
g19567 and n19527_not n19822_not ; n19823
g19568 and n19821_not n19823_not ; n19824
g19569 and n19821_not n19824_not ; n19825
g19570 and n19823_not n19824_not ; n19826
g19571 and n19825_not n19826_not ; n19827
g19572 and b[32] n8362 ; n19828
g19573 and b[30] n8715 ; n19829
g19574 and b[31] n8357 ; n19830
g19575 and n19829_not n19830_not ; n19831
g19576 and n19828_not n19831 ; n19832
g19577 and n4013 n8365 ; n19833
g19578 and n19832 n19833_not ; n19834
g19579 and a[50] n19834_not ; n19835
g19580 and a[50] n19835_not ; n19836
g19581 and n19834_not n19835_not ; n19837
g19582 and n19836_not n19837_not ; n19838
g19583 and n19827_not n19838 ; n19839
g19584 and n19827 n19838_not ; n19840
g19585 and n19839_not n19840_not ; n19841
g19586 and n19530_not n19533_not ; n19842
g19587 and n19841 n19842 ; n19843
g19588 and n19841_not n19842_not ; n19844
g19589 and n19843_not n19844_not ; n19845
g19590 and b[35] n7446 ; n19846
g19591 and b[33] n7787 ; n19847
g19592 and b[34] n7441 ; n19848
g19593 and n19847_not n19848_not ; n19849
g19594 and n19846_not n19849 ; n19850
g19595 and n4696 n7449 ; n19851
g19596 and n19850 n19851_not ; n19852
g19597 and a[47] n19852_not ; n19853
g19598 and a[47] n19853_not ; n19854
g19599 and n19852_not n19853_not ; n19855
g19600 and n19854_not n19855_not ; n19856
g19601 and n19845 n19856_not ; n19857
g19602 and n19845 n19857_not ; n19858
g19603 and n19856_not n19857_not ; n19859
g19604 and n19858_not n19859_not ; n19860
g19605 and n19539_not n19553_not ; n19861
g19606 and n19860_not n19861_not ; n19862
g19607 and n19860_not n19862_not ; n19863
g19608 and n19861_not n19862_not ; n19864
g19609 and n19863_not n19864_not ; n19865
g19610 and b[38] n6595 ; n19866
g19611 and b[36] n6902 ; n19867
g19612 and b[37] n6590 ; n19868
g19613 and n19867_not n19868_not ; n19869
g19614 and n19866_not n19869 ; n19870
g19615 and n5205 n6598 ; n19871
g19616 and n19870 n19871_not ; n19872
g19617 and a[44] n19872_not ; n19873
g19618 and a[44] n19873_not ; n19874
g19619 and n19872_not n19873_not ; n19875
g19620 and n19874_not n19875_not ; n19876
g19621 and n19865_not n19876 ; n19877
g19622 and n19865 n19876_not ; n19878
g19623 and n19877_not n19878_not ; n19879
g19624 and n19744_not n19879_not ; n19880
g19625 and n19744 n19879 ; n19881
g19626 and n19880_not n19881_not ; n19882
g19627 and n19743_not n19882 ; n19883
g19628 and n19743 n19882_not ; n19884
g19629 and n19883_not n19884_not ; n19885
g19630 and n19732_not n19885 ; n19886
g19631 and n19732 n19885_not ; n19887
g19632 and n19886_not n19887_not ; n19888
g19633 and n19731_not n19888 ; n19889
g19634 and n19731 n19888_not ; n19890
g19635 and n19889_not n19890_not ; n19891
g19636 and n19720_not n19891 ; n19892
g19637 and n19720 n19891_not ; n19893
g19638 and n19892_not n19893_not ; n19894
g19639 and b[47] n4287 ; n19895
g19640 and b[45] n4532 ; n19896
g19641 and b[46] n4282 ; n19897
g19642 and n19896_not n19897_not ; n19898
g19643 and n19895_not n19898 ; n19899
g19644 and n4290 n7703 ; n19900
g19645 and n19899 n19900_not ; n19901
g19646 and a[35] n19901_not ; n19902
g19647 and a[35] n19902_not ; n19903
g19648 and n19901_not n19902_not ; n19904
g19649 and n19903_not n19904_not ; n19905
g19650 and n19894 n19905_not ; n19906
g19651 and n19894 n19906_not ; n19907
g19652 and n19905_not n19906_not ; n19908
g19653 and n19907_not n19908_not ; n19909
g19654 and n19719 n19909_not ; n19910
g19655 and n19719_not n19909 ; n19911
g19656 and n19704_not n19911_not ; n19912
g19657 and n19910_not n19912 ; n19913
g19658 and n19704_not n19913_not ; n19914
g19659 and n19911_not n19913_not ; n19915
g19660 and n19910_not n19915 ; n19916
g19661 and n19914_not n19916_not ; n19917
g19662 and n19688 n19917_not ; n19918
g19663 and n19688_not n19917 ; n19919
g19664 and n19673_not n19919_not ; n19920
g19665 and n19918_not n19920 ; n19921
g19666 and n19673_not n19921_not ; n19922
g19667 and n19919_not n19921_not ; n19923
g19668 and n19918_not n19923 ; n19924
g19669 and n19922_not n19924_not ; n19925
g19670 and n19657_not n19925 ; n19926
g19671 and n19657 n19925_not ; n19927
g19672 and n19926_not n19927_not ; n19928
g19673 and n19642_not n19928 ; n19929
g19674 and n19642 n19928_not ; n19930
g19675 and n19929_not n19930_not ; n19931
g19676 and n19630_not n19931 ; n19932
g19677 and n19630_not n19932_not ; n19933
g19678 and n19931 n19932_not ; n19934
g19679 and n19933_not n19934_not ; n19935
g19680 and n19629_not n19935_not ; n19936
g19681 and n19629 n19934_not ; n19937
g19682 and n19933_not n19937 ; n19938
g19683 and n19936_not n19938_not ; f[80]
g19684 and n19932_not n19936_not ; n19940
g19685 and n19639_not n19929_not ; n19941
g19686 and n19656_not n19927_not ; n19942
g19687 and b[63] n1627 ; n19943
g19688 and b[61] n1763 ; n19944
g19689 and b[62] n1622 ; n19945
g19690 and n19944_not n19945_not ; n19946
g19691 and n19943_not n19946 ; n19947
g19692 and n1630 n13771 ; n19948
g19693 and n19947 n19948_not ; n19949
g19694 and a[20] n19949_not ; n19950
g19695 and a[20] n19950_not ; n19951
g19696 and n19949_not n19950_not ; n19952
g19697 and n19951_not n19952_not ; n19953
g19698 and n19942_not n19953_not ; n19954
g19699 and n19942_not n19954_not ; n19955
g19700 and n19953_not n19954_not ; n19956
g19701 and n19955_not n19956_not ; n19957
g19702 and b[60] n2048 ; n19958
g19703 and b[58] n2198 ; n19959
g19704 and b[59] n2043 ; n19960
g19705 and n19959_not n19960_not ; n19961
g19706 and n19958_not n19961 ; n19962
g19707 and n2051 n12211 ; n19963
g19708 and n19962 n19963_not ; n19964
g19709 and a[23] n19964_not ; n19965
g19710 and a[23] n19965_not ; n19966
g19711 and n19964_not n19965_not ; n19967
g19712 and n19966_not n19967_not ; n19968
g19713 and n19670_not n19921_not ; n19969
g19714 and n19968 n19969 ; n19970
g19715 and n19968_not n19969_not ; n19971
g19716 and n19970_not n19971_not ; n19972
g19717 and b[54] n3050 ; n19973
g19718 and b[52] n3243 ; n19974
g19719 and b[53] n3045 ; n19975
g19720 and n19974_not n19975_not ; n19976
g19721 and n19973_not n19976 ; n19977
g19722 and n3053 n9998 ; n19978
g19723 and n19977 n19978_not ; n19979
g19724 and a[29] n19979_not ; n19980
g19725 and a[29] n19980_not ; n19981
g19726 and n19979_not n19980_not ; n19982
g19727 and n19981_not n19982_not ; n19983
g19728 and n19701_not n19913_not ; n19984
g19729 and n19983 n19984 ; n19985
g19730 and n19983_not n19984_not ; n19986
g19731 and n19985_not n19986_not ; n19987
g19732 and n19880_not n19883_not ; n19988
g19733 and n19865_not n19876_not ; n19989
g19734 and n19862_not n19989_not ; n19990
g19735 and n19844_not n19857_not ; n19991
g19736 and b[27] n10426 ; n19992
g19737 and b[25] n10796 ; n19993
g19738 and b[26] n10421 ; n19994
g19739 and n19993_not n19994_not ; n19995
g19740 and n19992_not n19995 ; n19996
g19741 and n2990 n10429 ; n19997
g19742 and n19996 n19997_not ; n19998
g19743 and a[56] n19998_not ; n19999
g19744 and a[56] n19999_not ; n20000
g19745 and n19998_not n19999_not ; n20001
g19746 and n20000_not n20001_not ; n20002
g19747 and n19782_not n19796_not ; n20003
g19748 and b[21] n12668 ; n20004
g19749 and b[19] n13047 ; n20005
g19750 and b[20] n12663 ; n20006
g19751 and n20005_not n20006_not ; n20007
g19752 and n20004_not n20007 ; n20008
g19753 and n1984 n12671 ; n20009
g19754 and n20008 n20009_not ; n20010
g19755 and a[62] n20010_not ; n20011
g19756 and a[62] n20011_not ; n20012
g19757 and n20010_not n20011_not ; n20013
g19758 and n20012_not n20013_not ; n20014
g19759 and b[17] n13903 ; n20015
g19760 and b[18] n13488_not ; n20016
g19761 and n20015_not n20016_not ; n20017
g19762 and a[17]_not n20017_not ; n20018
g19763 and a[17] n20017 ; n20019
g19764 and n20018_not n20019_not ; n20020
g19765 and n19771_not n20020 ; n20021
g19766 and n19771 n20020_not ; n20022
g19767 and n20021_not n20022_not ; n20023
g19768 and n20014_not n20023 ; n20024
g19769 and n20014_not n20024_not ; n20025
g19770 and n20023 n20024_not ; n20026
g19771 and n20025_not n20026_not ; n20027
g19772 and n19777_not n20027_not ; n20028
g19773 and n19777_not n20028_not ; n20029
g19774 and n20027_not n20028_not ; n20030
g19775 and n20029_not n20030_not ; n20031
g19776 and b[24] n11531 ; n20032
g19777 and b[22] n11896 ; n20033
g19778 and b[23] n11526 ; n20034
g19779 and n20033_not n20034_not ; n20035
g19780 and n20032_not n20035 ; n20036
g19781 and n2458 n11534 ; n20037
g19782 and n20036 n20037_not ; n20038
g19783 and a[59] n20038_not ; n20039
g19784 and a[59] n20039_not ; n20040
g19785 and n20038_not n20039_not ; n20041
g19786 and n20040_not n20041_not ; n20042
g19787 and n20031 n20042 ; n20043
g19788 and n20031_not n20042_not ; n20044
g19789 and n20043_not n20044_not ; n20045
g19790 and n20003_not n20045 ; n20046
g19791 and n20003 n20045_not ; n20047
g19792 and n20046_not n20047_not ; n20048
g19793 and n20002_not n20048 ; n20049
g19794 and n20048 n20049_not ; n20050
g19795 and n20002_not n20049_not ; n20051
g19796 and n20050_not n20051_not ; n20052
g19797 and n19798_not n19801_not ; n20053
g19798 and n20052 n20053 ; n20054
g19799 and n20052_not n20053_not ; n20055
g19800 and n20054_not n20055_not ; n20056
g19801 and b[30] n9339 ; n20057
g19802 and b[28] n9732 ; n20058
g19803 and b[29] n9334 ; n20059
g19804 and n20058_not n20059_not ; n20060
g19805 and n20057_not n20060 ; n20061
g19806 and n3577 n9342 ; n20062
g19807 and n20061 n20062_not ; n20063
g19808 and a[53] n20063_not ; n20064
g19809 and a[53] n20064_not ; n20065
g19810 and n20063_not n20064_not ; n20066
g19811 and n20065_not n20066_not ; n20067
g19812 and n20056 n20067_not ; n20068
g19813 and n20056 n20068_not ; n20069
g19814 and n20067_not n20068_not ; n20070
g19815 and n20069_not n20070_not ; n20071
g19816 and n19804_not n19818_not ; n20072
g19817 and n20071 n20072 ; n20073
g19818 and n20071_not n20072_not ; n20074
g19819 and n20073_not n20074_not ; n20075
g19820 and b[33] n8362 ; n20076
g19821 and b[31] n8715 ; n20077
g19822 and b[32] n8357 ; n20078
g19823 and n20077_not n20078_not ; n20079
g19824 and n20076_not n20079 ; n20080
g19825 and n4223 n8365 ; n20081
g19826 and n20080 n20081_not ; n20082
g19827 and a[50] n20082_not ; n20083
g19828 and a[50] n20083_not ; n20084
g19829 and n20082_not n20083_not ; n20085
g19830 and n20084_not n20085_not ; n20086
g19831 and n19827_not n19838_not ; n20087
g19832 and n19824_not n20087_not ; n20088
g19833 and n20086_not n20088_not ; n20089
g19834 and n20086 n20088 ; n20090
g19835 and n20089_not n20090_not ; n20091
g19836 and n20075_not n20091 ; n20092
g19837 and n20075 n20091_not ; n20093
g19838 and n20092_not n20093_not ; n20094
g19839 and b[36] n7446 ; n20095
g19840 and b[34] n7787 ; n20096
g19841 and b[35] n7441 ; n20097
g19842 and n20096_not n20097_not ; n20098
g19843 and n20095_not n20098 ; n20099
g19844 and n4922 n7449 ; n20100
g19845 and n20099 n20100_not ; n20101
g19846 and a[47] n20101_not ; n20102
g19847 and a[47] n20102_not ; n20103
g19848 and n20101_not n20102_not ; n20104
g19849 and n20103_not n20104_not ; n20105
g19850 and n20094_not n20105_not ; n20106
g19851 and n20094 n20105 ; n20107
g19852 and n20106_not n20107_not ; n20108
g19853 and n19991 n20108_not ; n20109
g19854 and n19991_not n20108 ; n20110
g19855 and n20109_not n20110_not ; n20111
g19856 and b[39] n6595 ; n20112
g19857 and b[37] n6902 ; n20113
g19858 and b[38] n6590 ; n20114
g19859 and n20113_not n20114_not ; n20115
g19860 and n20112_not n20115 ; n20116
g19861 and n5451 n6598 ; n20117
g19862 and n20116 n20117_not ; n20118
g19863 and a[44] n20118_not ; n20119
g19864 and a[44] n20119_not ; n20120
g19865 and n20118_not n20119_not ; n20121
g19866 and n20120_not n20121_not ; n20122
g19867 and n20111 n20122_not ; n20123
g19868 and n20111 n20123_not ; n20124
g19869 and n20122_not n20123_not ; n20125
g19870 and n20124_not n20125_not ; n20126
g19871 and n19990_not n20126 ; n20127
g19872 and n19990 n20126_not ; n20128
g19873 and n20127_not n20128_not ; n20129
g19874 and b[42] n5777 ; n20130
g19875 and b[40] n6059 ; n20131
g19876 and b[41] n5772 ; n20132
g19877 and n20131_not n20132_not ; n20133
g19878 and n20130_not n20133 ; n20134
g19879 and n5780 n6489 ; n20135
g19880 and n20134 n20135_not ; n20136
g19881 and a[41] n20136_not ; n20137
g19882 and a[41] n20137_not ; n20138
g19883 and n20136_not n20137_not ; n20139
g19884 and n20138_not n20139_not ; n20140
g19885 and n20129_not n20140_not ; n20141
g19886 and n20129 n20140 ; n20142
g19887 and n20141_not n20142_not ; n20143
g19888 and n19988 n20143_not ; n20144
g19889 and n19988_not n20143 ; n20145
g19890 and n20144_not n20145_not ; n20146
g19891 and b[45] n5035 ; n20147
g19892 and b[43] n5277 ; n20148
g19893 and b[44] n5030 ; n20149
g19894 and n20148_not n20149_not ; n20150
g19895 and n20147_not n20150 ; n20151
g19896 and n5038 n7361 ; n20152
g19897 and n20151 n20152_not ; n20153
g19898 and a[38] n20153_not ; n20154
g19899 and a[38] n20154_not ; n20155
g19900 and n20153_not n20154_not ; n20156
g19901 and n20155_not n20156_not ; n20157
g19902 and n20146 n20157_not ; n20158
g19903 and n20146 n20158_not ; n20159
g19904 and n20157_not n20158_not ; n20160
g19905 and n20159_not n20160_not ; n20161
g19906 and n19886_not n19889_not ; n20162
g19907 and n20161 n20162 ; n20163
g19908 and n20161_not n20162_not ; n20164
g19909 and n20163_not n20164_not ; n20165
g19910 and b[48] n4287 ; n20166
g19911 and b[46] n4532 ; n20167
g19912 and b[47] n4282 ; n20168
g19913 and n20167_not n20168_not ; n20169
g19914 and n20166_not n20169 ; n20170
g19915 and n4290 n8009 ; n20171
g19916 and n20170 n20171_not ; n20172
g19917 and a[35] n20172_not ; n20173
g19918 and a[35] n20173_not ; n20174
g19919 and n20172_not n20173_not ; n20175
g19920 and n20174_not n20175_not ; n20176
g19921 and n20165 n20176_not ; n20177
g19922 and n20165 n20177_not ; n20178
g19923 and n20176_not n20177_not ; n20179
g19924 and n20178_not n20179_not ; n20180
g19925 and n19892_not n19906_not ; n20181
g19926 and n20180 n20181 ; n20182
g19927 and n20180_not n20181_not ; n20183
g19928 and n20182_not n20183_not ; n20184
g19929 and b[51] n3638 ; n20185
g19930 and b[49] n3843 ; n20186
g19931 and b[50] n3633 ; n20187
g19932 and n20186_not n20187_not ; n20188
g19933 and n20185_not n20188 ; n20189
g19934 and n3641 n8976 ; n20190
g19935 and n20189 n20190_not ; n20191
g19936 and a[32] n20191_not ; n20192
g19937 and a[32] n20192_not ; n20193
g19938 and n20191_not n20192_not ; n20194
g19939 and n20193_not n20194_not ; n20195
g19940 and n19718_not n19910_not ; n20196
g19941 and n20195_not n20196_not ; n20197
g19942 and n20195 n20196 ; n20198
g19943 and n20197_not n20198_not ; n20199
g19944 and n20184 n20199 ; n20200
g19945 and n20184 n20200_not ; n20201
g19946 and n20199 n20200_not ; n20202
g19947 and n20201_not n20202_not ; n20203
g19948 and n19987 n20203_not ; n20204
g19949 and n19987 n20204_not ; n20205
g19950 and n20203_not n20204_not ; n20206
g19951 and n20205_not n20206_not ; n20207
g19952 and b[57] n2539 ; n20208
g19953 and b[55] n2685 ; n20209
g19954 and b[56] n2534 ; n20210
g19955 and n20209_not n20210_not ; n20211
g19956 and n20208_not n20211 ; n20212
g19957 and n2542 n11410 ; n20213
g19958 and n20212 n20213_not ; n20214
g19959 and a[26] n20214_not ; n20215
g19960 and a[26] n20215_not ; n20216
g19961 and n20214_not n20215_not ; n20217
g19962 and n20216_not n20217_not ; n20218
g19963 and n19687_not n19918_not ; n20219
g19964 and n20218_not n20219_not ; n20220
g19965 and n20218 n20219 ; n20221
g19966 and n20220_not n20221_not ; n20222
g19967 and n20207_not n20222 ; n20223
g19968 and n20207_not n20223_not ; n20224
g19969 and n20222 n20223_not ; n20225
g19970 and n20224_not n20225_not ; n20226
g19971 and n19972 n20226_not ; n20227
g19972 and n19972 n20227_not ; n20228
g19973 and n20226_not n20227_not ; n20229
g19974 and n20228_not n20229_not ; n20230
g19975 and n19957_not n20230 ; n20231
g19976 and n19957 n20230_not ; n20232
g19977 and n20231_not n20232_not ; n20233
g19978 and n19941_not n20233_not ; n20234
g19979 and n19941_not n20234_not ; n20235
g19980 and n20233_not n20234_not ; n20236
g19981 and n20235_not n20236_not ; n20237
g19982 and n19940_not n20237_not ; n20238
g19983 and n19940 n20236_not ; n20239
g19984 and n20235_not n20239 ; n20240
g19985 and n20238_not n20240_not ; f[81]
g19986 and n20234_not n20238_not ; n20242
g19987 and n19957_not n20230_not ; n20243
g19988 and n19954_not n20243_not ; n20244
g19989 and b[61] n2048 ; n20245
g19990 and b[59] n2198 ; n20246
g19991 and b[60] n2043 ; n20247
g19992 and n20246_not n20247_not ; n20248
g19993 and n20245_not n20248 ; n20249
g19994 and n2051 n12969 ; n20250
g19995 and n20249 n20250_not ; n20251
g19996 and a[23] n20251_not ; n20252
g19997 and a[23] n20252_not ; n20253
g19998 and n20251_not n20252_not ; n20254
g19999 and n20253_not n20254_not ; n20255
g20000 and n20220_not n20223_not ; n20256
g20001 and n20255 n20256 ; n20257
g20002 and n20255_not n20256_not ; n20258
g20003 and n20257_not n20258_not ; n20259
g20004 and b[58] n2539 ; n20260
g20005 and b[56] n2685 ; n20261
g20006 and b[57] n2534 ; n20262
g20007 and n20261_not n20262_not ; n20263
g20008 and n20260_not n20263 ; n20264
g20009 and n2542 n11436 ; n20265
g20010 and n20264 n20265_not ; n20266
g20011 and a[26] n20266_not ; n20267
g20012 and a[26] n20267_not ; n20268
g20013 and n20266_not n20267_not ; n20269
g20014 and n20268_not n20269_not ; n20270
g20015 and n19986_not n20204_not ; n20271
g20016 and n20270 n20271 ; n20272
g20017 and n20270_not n20271_not ; n20273
g20018 and n20272_not n20273_not ; n20274
g20019 and b[55] n3050 ; n20275
g20020 and b[53] n3243 ; n20276
g20021 and b[54] n3045 ; n20277
g20022 and n20276_not n20277_not ; n20278
g20023 and n20275_not n20278 ; n20279
g20024 and n3053 n10684 ; n20280
g20025 and n20279 n20280_not ; n20281
g20026 and a[29] n20281_not ; n20282
g20027 and a[29] n20282_not ; n20283
g20028 and n20281_not n20282_not ; n20284
g20029 and n20283_not n20284_not ; n20285
g20030 and n20197_not n20200_not ; n20286
g20031 and n20285 n20286 ; n20287
g20032 and n20285_not n20286_not ; n20288
g20033 and n20287_not n20288_not ; n20289
g20034 and b[52] n3638 ; n20290
g20035 and b[50] n3843 ; n20291
g20036 and b[51] n3633 ; n20292
g20037 and n20291_not n20292_not ; n20293
g20038 and n20290_not n20293 ; n20294
g20039 and n3641 n9628 ; n20295
g20040 and n20294 n20295_not ; n20296
g20041 and a[32] n20296_not ; n20297
g20042 and a[32] n20297_not ; n20298
g20043 and n20296_not n20297_not ; n20299
g20044 and n20298_not n20299_not ; n20300
g20045 and n20177_not n20183_not ; n20301
g20046 and n20300 n20301 ; n20302
g20047 and n20300_not n20301_not ; n20303
g20048 and n20302_not n20303_not ; n20304
g20049 and b[43] n5777 ; n20305
g20050 and b[41] n6059 ; n20306
g20051 and b[42] n5772 ; n20307
g20052 and n20306_not n20307_not ; n20308
g20053 and n20305_not n20308 ; n20309
g20054 and n5780 n6515 ; n20310
g20055 and n20309 n20310_not ; n20311
g20056 and a[41] n20311_not ; n20312
g20057 and a[41] n20312_not ; n20313
g20058 and n20311_not n20312_not ; n20314
g20059 and n20313_not n20314_not ; n20315
g20060 and n19990_not n20126_not ; n20316
g20061 and n20123_not n20316_not ; n20317
g20062 and b[40] n6595 ; n20318
g20063 and b[38] n6902 ; n20319
g20064 and b[39] n6590 ; n20320
g20065 and n20319_not n20320_not ; n20321
g20066 and n20318_not n20321 ; n20322
g20067 and n5955 n6598 ; n20323
g20068 and n20322 n20323_not ; n20324
g20069 and a[44] n20324_not ; n20325
g20070 and a[44] n20325_not ; n20326
g20071 and n20324_not n20325_not ; n20327
g20072 and n20326_not n20327_not ; n20328
g20073 and n20106_not n20110_not ; n20329
g20074 and b[31] n9339 ; n20330
g20075 and b[29] n9732 ; n20331
g20076 and b[30] n9334 ; n20332
g20077 and n20331_not n20332_not ; n20333
g20078 and n20330_not n20333 ; n20334
g20079 and n3796 n9342 ; n20335
g20080 and n20334 n20335_not ; n20336
g20081 and a[53] n20336_not ; n20337
g20082 and a[53] n20337_not ; n20338
g20083 and n20336_not n20337_not ; n20339
g20084 and n20338_not n20339_not ; n20340
g20085 and n20044_not n20046_not ; n20341
g20086 and b[25] n11531 ; n20342
g20087 and b[23] n11896 ; n20343
g20088 and b[24] n11526 ; n20344
g20089 and n20343_not n20344_not ; n20345
g20090 and n20342_not n20345 ; n20346
g20091 and n2485 n11534 ; n20347
g20092 and n20346 n20347_not ; n20348
g20093 and a[59] n20348_not ; n20349
g20094 and a[59] n20349_not ; n20350
g20095 and n20348_not n20349_not ; n20351
g20096 and n20350_not n20351_not ; n20352
g20097 and b[18] n13903 ; n20353
g20098 and b[19] n13488_not ; n20354
g20099 and n20353_not n20354_not ; n20355
g20100 and n20018_not n20021_not ; n20356
g20101 and n20355_not n20356 ; n20357
g20102 and n20355 n20356_not ; n20358
g20103 and n20357_not n20358_not ; n20359
g20104 and b[22] n12668 ; n20360
g20105 and b[20] n13047 ; n20361
g20106 and b[21] n12663 ; n20362
g20107 and n20361_not n20362_not ; n20363
g20108 and n20360_not n20363 ; n20364
g20109 and n2145 n12671 ; n20365
g20110 and n20364 n20365_not ; n20366
g20111 and a[62] n20366_not ; n20367
g20112 and a[62] n20367_not ; n20368
g20113 and n20366_not n20367_not ; n20369
g20114 and n20368_not n20369_not ; n20370
g20115 and n20359_not n20370 ; n20371
g20116 and n20359 n20370_not ; n20372
g20117 and n20371_not n20372_not ; n20373
g20118 and n20024_not n20028_not ; n20374
g20119 and n20373 n20374_not ; n20375
g20120 and n20373_not n20374 ; n20376
g20121 and n20375_not n20376_not ; n20377
g20122 and n20352_not n20377 ; n20378
g20123 and n20377 n20378_not ; n20379
g20124 and n20352_not n20378_not ; n20380
g20125 and n20379_not n20380_not ; n20381
g20126 and n20341_not n20381 ; n20382
g20127 and n20341 n20381_not ; n20383
g20128 and n20382_not n20383_not ; n20384
g20129 and b[28] n10426 ; n20385
g20130 and b[26] n10796 ; n20386
g20131 and b[27] n10421 ; n20387
g20132 and n20386_not n20387_not ; n20388
g20133 and n20385_not n20388 ; n20389
g20134 and n3189 n10429 ; n20390
g20135 and n20389 n20390_not ; n20391
g20136 and a[56] n20391_not ; n20392
g20137 and a[56] n20392_not ; n20393
g20138 and n20391_not n20392_not ; n20394
g20139 and n20393_not n20394_not ; n20395
g20140 and n20384 n20395 ; n20396
g20141 and n20384_not n20395_not ; n20397
g20142 and n20396_not n20397_not ; n20398
g20143 and n20049_not n20055_not ; n20399
g20144 and n20398 n20399_not ; n20400
g20145 and n20398_not n20399 ; n20401
g20146 and n20400_not n20401_not ; n20402
g20147 and n20340_not n20402 ; n20403
g20148 and n20402 n20403_not ; n20404
g20149 and n20340_not n20403_not ; n20405
g20150 and n20404_not n20405_not ; n20406
g20151 and n20068_not n20074_not ; n20407
g20152 and n20406 n20407 ; n20408
g20153 and n20406_not n20407_not ; n20409
g20154 and n20408_not n20409_not ; n20410
g20155 and b[34] n8362 ; n20411
g20156 and b[32] n8715 ; n20412
g20157 and b[33] n8357 ; n20413
g20158 and n20412_not n20413_not ; n20414
g20159 and n20411_not n20414 ; n20415
g20160 and n4466 n8365 ; n20416
g20161 and n20415 n20416_not ; n20417
g20162 and a[50] n20417_not ; n20418
g20163 and a[50] n20418_not ; n20419
g20164 and n20417_not n20418_not ; n20420
g20165 and n20419_not n20420_not ; n20421
g20166 and n20410 n20421_not ; n20422
g20167 and n20410 n20422_not ; n20423
g20168 and n20421_not n20422_not ; n20424
g20169 and n20423_not n20424_not ; n20425
g20170 and n20075 n20091 ; n20426
g20171 and n20089_not n20426_not ; n20427
g20172 and n20425 n20427 ; n20428
g20173 and n20425_not n20427_not ; n20429
g20174 and n20428_not n20429_not ; n20430
g20175 and b[37] n7446 ; n20431
g20176 and b[35] n7787 ; n20432
g20177 and b[36] n7441 ; n20433
g20178 and n20432_not n20433_not ; n20434
g20179 and n20431_not n20434 ; n20435
g20180 and n5181 n7449 ; n20436
g20181 and n20435 n20436_not ; n20437
g20182 and a[47] n20437_not ; n20438
g20183 and a[47] n20438_not ; n20439
g20184 and n20437_not n20438_not ; n20440
g20185 and n20439_not n20440_not ; n20441
g20186 and n20430_not n20441 ; n20442
g20187 and n20430 n20441_not ; n20443
g20188 and n20442_not n20443_not ; n20444
g20189 and n20329_not n20444 ; n20445
g20190 and n20329_not n20445_not ; n20446
g20191 and n20444 n20445_not ; n20447
g20192 and n20446_not n20447_not ; n20448
g20193 and n20328_not n20448_not ; n20449
g20194 and n20328 n20447_not ; n20450
g20195 and n20446_not n20450 ; n20451
g20196 and n20449_not n20451_not ; n20452
g20197 and n20317_not n20452 ; n20453
g20198 and n20317 n20452_not ; n20454
g20199 and n20453_not n20454_not ; n20455
g20200 and n20315_not n20455 ; n20456
g20201 and n20455 n20456_not ; n20457
g20202 and n20315_not n20456_not ; n20458
g20203 and n20457_not n20458_not ; n20459
g20204 and n20141_not n20145_not ; n20460
g20205 and n20459 n20460 ; n20461
g20206 and n20459_not n20460_not ; n20462
g20207 and n20461_not n20462_not ; n20463
g20208 and b[46] n5035 ; n20464
g20209 and b[44] n5277 ; n20465
g20210 and b[45] n5030 ; n20466
g20211 and n20465_not n20466_not ; n20467
g20212 and n20464_not n20467 ; n20468
g20213 and n5038 n7677 ; n20469
g20214 and n20468 n20469_not ; n20470
g20215 and a[38] n20470_not ; n20471
g20216 and a[38] n20471_not ; n20472
g20217 and n20470_not n20471_not ; n20473
g20218 and n20472_not n20473_not ; n20474
g20219 and n20463 n20474_not ; n20475
g20220 and n20463 n20475_not ; n20476
g20221 and n20474_not n20475_not ; n20477
g20222 and n20476_not n20477_not ; n20478
g20223 and n20158_not n20164_not ; n20479
g20224 and n20478 n20479 ; n20480
g20225 and n20478_not n20479_not ; n20481
g20226 and n20480_not n20481_not ; n20482
g20227 and b[49] n4287 ; n20483
g20228 and b[47] n4532 ; n20484
g20229 and b[48] n4282 ; n20485
g20230 and n20484_not n20485_not ; n20486
g20231 and n20483_not n20486 ; n20487
g20232 and n4290 n8625 ; n20488
g20233 and n20487 n20488_not ; n20489
g20234 and a[35] n20489_not ; n20490
g20235 and a[35] n20490_not ; n20491
g20236 and n20489_not n20490_not ; n20492
g20237 and n20491_not n20492_not ; n20493
g20238 and n20482 n20493_not ; n20494
g20239 and n20482 n20494_not ; n20495
g20240 and n20493_not n20494_not ; n20496
g20241 and n20495_not n20496_not ; n20497
g20242 and n20304 n20497_not ; n20498
g20243 and n20304_not n20497 ; n20499
g20244 and n20289 n20499_not ; n20500
g20245 and n20498_not n20500 ; n20501
g20246 and n20289 n20501_not ; n20502
g20247 and n20499_not n20501_not ; n20503
g20248 and n20498_not n20503 ; n20504
g20249 and n20502_not n20504_not ; n20505
g20250 and n20274 n20505_not ; n20506
g20251 and n20274_not n20505 ; n20507
g20252 and n20259 n20507_not ; n20508
g20253 and n20506_not n20508 ; n20509
g20254 and n20259 n20509_not ; n20510
g20255 and n20507_not n20509_not ; n20511
g20256 and n20506_not n20511 ; n20512
g20257 and n20510_not n20512_not ; n20513
g20258 and n19971_not n20227_not ; n20514
g20259 and b[62] n1763 ; n20515
g20260 and b[63] n1622 ; n20516
g20261 and n20515_not n20516_not ; n20517
g20262 and n1630_not n20517 ; n20518
g20263 and n13800 n20517 ; n20519
g20264 and n20518_not n20519_not ; n20520
g20265 and a[20] n20520_not ; n20521
g20266 and a[20]_not n20520 ; n20522
g20267 and n20521_not n20522_not ; n20523
g20268 and n20514_not n20523_not ; n20524
g20269 and n20514_not n20524_not ; n20525
g20270 and n20523_not n20524_not ; n20526
g20271 and n20525_not n20526_not ; n20527
g20272 and n20513_not n20527_not ; n20528
g20273 and n20513 n20526_not ; n20529
g20274 and n20525_not n20529 ; n20530
g20275 and n20528_not n20530_not ; n20531
g20276 and n20244_not n20531 ; n20532
g20277 and n20244_not n20532_not ; n20533
g20278 and n20531 n20532_not ; n20534
g20279 and n20533_not n20534_not ; n20535
g20280 and n20242_not n20535_not ; n20536
g20281 and n20242 n20534_not ; n20537
g20282 and n20533_not n20537 ; n20538
g20283 and n20536_not n20538_not ; f[82]
g20284 and n20532_not n20536_not ; n20540
g20285 and n20524_not n20528_not ; n20541
g20286 and n20258_not n20509_not ; n20542
g20287 and b[63] n1763 ; n20543
g20288 and n1630 n13797 ; n20544
g20289 and n20543_not n20544_not ; n20545
g20290 and a[20] n20545_not ; n20546
g20291 and a[20] n20546_not ; n20547
g20292 and n20545_not n20546_not ; n20548
g20293 and n20547_not n20548_not ; n20549
g20294 and n20542_not n20549_not ; n20550
g20295 and n20542_not n20550_not ; n20551
g20296 and n20549_not n20550_not ; n20552
g20297 and n20551_not n20552_not ; n20553
g20298 and b[62] n2048 ; n20554
g20299 and b[60] n2198 ; n20555
g20300 and b[61] n2043 ; n20556
g20301 and n20555_not n20556_not ; n20557
g20302 and n20554_not n20557 ; n20558
g20303 and n2051 n13370 ; n20559
g20304 and n20558 n20559_not ; n20560
g20305 and a[23] n20560_not ; n20561
g20306 and a[23] n20561_not ; n20562
g20307 and n20560_not n20561_not ; n20563
g20308 and n20562_not n20563_not ; n20564
g20309 and n20273_not n20506_not ; n20565
g20310 and n20564_not n20565_not ; n20566
g20311 and n20564_not n20566_not ; n20567
g20312 and n20565_not n20566_not ; n20568
g20313 and n20567_not n20568_not ; n20569
g20314 and b[59] n2539 ; n20570
g20315 and b[57] n2685 ; n20571
g20316 and b[58] n2534 ; n20572
g20317 and n20571_not n20572_not ; n20573
g20318 and n20570_not n20573 ; n20574
g20319 and n2542 n12179 ; n20575
g20320 and n20574 n20575_not ; n20576
g20321 and a[26] n20576_not ; n20577
g20322 and a[26] n20577_not ; n20578
g20323 and n20576_not n20577_not ; n20579
g20324 and n20578_not n20579_not ; n20580
g20325 and n20288_not n20501_not ; n20581
g20326 and n20580 n20581 ; n20582
g20327 and n20580_not n20581_not ; n20583
g20328 and n20582_not n20583_not ; n20584
g20329 and b[56] n3050 ; n20585
g20330 and b[54] n3243 ; n20586
g20331 and b[55] n3045 ; n20587
g20332 and n20586_not n20587_not ; n20588
g20333 and n20585_not n20588 ; n20589
g20334 and n3053 n10708 ; n20590
g20335 and n20589 n20590_not ; n20591
g20336 and a[29] n20591_not ; n20592
g20337 and a[29] n20592_not ; n20593
g20338 and n20591_not n20592_not ; n20594
g20339 and n20593_not n20594_not ; n20595
g20340 and n20303_not n20498_not ; n20596
g20341 and n20595_not n20596_not ; n20597
g20342 and n20595_not n20597_not ; n20598
g20343 and n20596_not n20597_not ; n20599
g20344 and n20598_not n20599_not ; n20600
g20345 and b[53] n3638 ; n20601
g20346 and b[51] n3843 ; n20602
g20347 and b[52] n3633 ; n20603
g20348 and n20602_not n20603_not ; n20604
g20349 and n20601_not n20604 ; n20605
g20350 and n3641 n9972 ; n20606
g20351 and n20605 n20606_not ; n20607
g20352 and a[32] n20607_not ; n20608
g20353 and a[32] n20608_not ; n20609
g20354 and n20607_not n20608_not ; n20610
g20355 and n20609_not n20610_not ; n20611
g20356 and n20481_not n20494_not ; n20612
g20357 and n20611 n20612 ; n20613
g20358 and n20611_not n20612_not ; n20614
g20359 and n20613_not n20614_not ; n20615
g20360 and n20453_not n20456_not ; n20616
g20361 and b[44] n5777 ; n20617
g20362 and b[42] n6059 ; n20618
g20363 and b[43] n5772 ; n20619
g20364 and n20618_not n20619_not ; n20620
g20365 and n20617_not n20620 ; n20621
g20366 and n5780 n7072 ; n20622
g20367 and n20621 n20622_not ; n20623
g20368 and a[41] n20623_not ; n20624
g20369 and a[41] n20624_not ; n20625
g20370 and n20623_not n20624_not ; n20626
g20371 and n20625_not n20626_not ; n20627
g20372 and n20445_not n20449_not ; n20628
g20373 and b[41] n6595 ; n20629
g20374 and b[39] n6902 ; n20630
g20375 and b[40] n6590 ; n20631
g20376 and n20630_not n20631_not ; n20632
g20377 and n20629_not n20632 ; n20633
g20378 and n6219 n6598 ; n20634
g20379 and n20633 n20634_not ; n20635
g20380 and a[44] n20635_not ; n20636
g20381 and a[44] n20636_not ; n20637
g20382 and n20635_not n20636_not ; n20638
g20383 and n20637_not n20638_not ; n20639
g20384 and n20429_not n20443_not ; n20640
g20385 and b[38] n7446 ; n20641
g20386 and b[36] n7787 ; n20642
g20387 and b[37] n7441 ; n20643
g20388 and n20642_not n20643_not ; n20644
g20389 and n20641_not n20644 ; n20645
g20390 and n5205 n7449 ; n20646
g20391 and n20645 n20646_not ; n20647
g20392 and a[47] n20647_not ; n20648
g20393 and a[47] n20648_not ; n20649
g20394 and n20647_not n20648_not ; n20650
g20395 and n20649_not n20650_not ; n20651
g20396 and n20409_not n20422_not ; n20652
g20397 and b[35] n8362 ; n20653
g20398 and b[33] n8715 ; n20654
g20399 and b[34] n8357 ; n20655
g20400 and n20654_not n20655_not ; n20656
g20401 and n20653_not n20656 ; n20657
g20402 and n4696 n8365 ; n20658
g20403 and n20657 n20658_not ; n20659
g20404 and a[50] n20659_not ; n20660
g20405 and a[50] n20660_not ; n20661
g20406 and n20659_not n20660_not ; n20662
g20407 and n20661_not n20662_not ; n20663
g20408 and n20400_not n20403_not ; n20664
g20409 and n20375_not n20378_not ; n20665
g20410 and b[26] n11531 ; n20666
g20411 and b[24] n11896 ; n20667
g20412 and b[25] n11526 ; n20668
g20413 and n20667_not n20668_not ; n20669
g20414 and n20666_not n20669 ; n20670
g20415 and n2813 n11534 ; n20671
g20416 and n20670 n20671_not ; n20672
g20417 and a[59] n20672_not ; n20673
g20418 and a[59] n20673_not ; n20674
g20419 and n20672_not n20673_not ; n20675
g20420 and n20674_not n20675_not ; n20676
g20421 and n20358_not n20372_not ; n20677
g20422 and b[19] n13903 ; n20678
g20423 and b[20] n13488_not ; n20679
g20424 and n20678_not n20679_not ; n20680
g20425 and n20355_not n20680 ; n20681
g20426 and n20355 n20680_not ; n20682
g20427 and n20681_not n20682_not ; n20683
g20428 and b[23] n12668 ; n20684
g20429 and b[21] n13047 ; n20685
g20430 and b[22] n12663 ; n20686
g20431 and n20685_not n20686_not ; n20687
g20432 and n20684_not n20687 ; n20688
g20433 and n12671_not n20688 ; n20689
g20434 and n2300_not n20688 ; n20690
g20435 and n20689_not n20690_not ; n20691
g20436 and a[62] n20691_not ; n20692
g20437 and a[62]_not n20691 ; n20693
g20438 and n20692_not n20693_not ; n20694
g20439 and n20683 n20694_not ; n20695
g20440 and n20683_not n20694 ; n20696
g20441 and n20695_not n20696_not ; n20697
g20442 and n20677_not n20697 ; n20698
g20443 and n20677 n20697_not ; n20699
g20444 and n20698_not n20699_not ; n20700
g20445 and n20676_not n20700 ; n20701
g20446 and n20676 n20700_not ; n20702
g20447 and n20701_not n20702_not ; n20703
g20448 and n20665_not n20703 ; n20704
g20449 and n20665 n20703_not ; n20705
g20450 and n20704_not n20705_not ; n20706
g20451 and b[29] n10426 ; n20707
g20452 and b[27] n10796 ; n20708
g20453 and b[28] n10421 ; n20709
g20454 and n20708_not n20709_not ; n20710
g20455 and n20707_not n20710 ; n20711
g20456 and n3383 n10429 ; n20712
g20457 and n20711 n20712_not ; n20713
g20458 and a[56] n20713_not ; n20714
g20459 and a[56] n20714_not ; n20715
g20460 and n20713_not n20714_not ; n20716
g20461 and n20715_not n20716_not ; n20717
g20462 and n20706 n20717_not ; n20718
g20463 and n20706 n20718_not ; n20719
g20464 and n20717_not n20718_not ; n20720
g20465 and n20719_not n20720_not ; n20721
g20466 and n20341_not n20381_not ; n20722
g20467 and n20397_not n20722_not ; n20723
g20468 and n20721_not n20723_not ; n20724
g20469 and n20721_not n20724_not ; n20725
g20470 and n20723_not n20724_not ; n20726
g20471 and n20725_not n20726_not ; n20727
g20472 and b[32] n9339 ; n20728
g20473 and b[30] n9732 ; n20729
g20474 and b[31] n9334 ; n20730
g20475 and n20729_not n20730_not ; n20731
g20476 and n20728_not n20731 ; n20732
g20477 and n4013 n9342 ; n20733
g20478 and n20732 n20733_not ; n20734
g20479 and a[53] n20734_not ; n20735
g20480 and a[53] n20735_not ; n20736
g20481 and n20734_not n20735_not ; n20737
g20482 and n20736_not n20737_not ; n20738
g20483 and n20727_not n20738 ; n20739
g20484 and n20727 n20738_not ; n20740
g20485 and n20739_not n20740_not ; n20741
g20486 and n20664_not n20741_not ; n20742
g20487 and n20664 n20741 ; n20743
g20488 and n20742_not n20743_not ; n20744
g20489 and n20663_not n20744 ; n20745
g20490 and n20663 n20744_not ; n20746
g20491 and n20745_not n20746_not ; n20747
g20492 and n20652_not n20747 ; n20748
g20493 and n20652 n20747_not ; n20749
g20494 and n20748_not n20749_not ; n20750
g20495 and n20651_not n20750 ; n20751
g20496 and n20651 n20750_not ; n20752
g20497 and n20751_not n20752_not ; n20753
g20498 and n20640_not n20753 ; n20754
g20499 and n20640 n20753_not ; n20755
g20500 and n20754_not n20755_not ; n20756
g20501 and n20639_not n20756 ; n20757
g20502 and n20639 n20756_not ; n20758
g20503 and n20757_not n20758_not ; n20759
g20504 and n20628_not n20759 ; n20760
g20505 and n20628 n20759_not ; n20761
g20506 and n20760_not n20761_not ; n20762
g20507 and n20627_not n20762 ; n20763
g20508 and n20627 n20762_not ; n20764
g20509 and n20763_not n20764_not ; n20765
g20510 and n20616_not n20765 ; n20766
g20511 and n20616 n20765_not ; n20767
g20512 and n20766_not n20767_not ; n20768
g20513 and b[47] n5035 ; n20769
g20514 and b[45] n5277 ; n20770
g20515 and b[46] n5030 ; n20771
g20516 and n20770_not n20771_not ; n20772
g20517 and n20769_not n20772 ; n20773
g20518 and n5038 n7703 ; n20774
g20519 and n20773 n20774_not ; n20775
g20520 and a[38] n20775_not ; n20776
g20521 and a[38] n20776_not ; n20777
g20522 and n20775_not n20776_not ; n20778
g20523 and n20777_not n20778_not ; n20779
g20524 and n20768 n20779_not ; n20780
g20525 and n20768 n20780_not ; n20781
g20526 and n20779_not n20780_not ; n20782
g20527 and n20781_not n20782_not ; n20783
g20528 and n20462_not n20475_not ; n20784
g20529 and n20783 n20784 ; n20785
g20530 and n20783_not n20784_not ; n20786
g20531 and n20785_not n20786_not ; n20787
g20532 and b[50] n4287 ; n20788
g20533 and b[48] n4532 ; n20789
g20534 and b[49] n4282 ; n20790
g20535 and n20789_not n20790_not ; n20791
g20536 and n20788_not n20791 ; n20792
g20537 and n4290 n8949 ; n20793
g20538 and n20792 n20793_not ; n20794
g20539 and a[35] n20794_not ; n20795
g20540 and a[35] n20795_not ; n20796
g20541 and n20794_not n20795_not ; n20797
g20542 and n20796_not n20797_not ; n20798
g20543 and n20787 n20798_not ; n20799
g20544 and n20787_not n20798 ; n20800
g20545 and n20615 n20800_not ; n20801
g20546 and n20799_not n20801 ; n20802
g20547 and n20615 n20802_not ; n20803
g20548 and n20800_not n20802_not ; n20804
g20549 and n20799_not n20804 ; n20805
g20550 and n20803_not n20805_not ; n20806
g20551 and n20600_not n20806 ; n20807
g20552 and n20600 n20806_not ; n20808
g20553 and n20807_not n20808_not ; n20809
g20554 and n20584 n20809_not ; n20810
g20555 and n20584 n20810_not ; n20811
g20556 and n20809_not n20810_not ; n20812
g20557 and n20811_not n20812_not ; n20813
g20558 and n20569_not n20813 ; n20814
g20559 and n20569 n20813_not ; n20815
g20560 and n20814_not n20815_not ; n20816
g20561 and n20553_not n20816_not ; n20817
g20562 and n20553 n20816 ; n20818
g20563 and n20817_not n20818_not ; n20819
g20564 and n20541_not n20819 ; n20820
g20565 and n20541 n20819_not ; n20821
g20566 and n20820_not n20821_not ; n20822
g20567 and n20540_not n20822 ; n20823
g20568 and n20540 n20822_not ; n20824
g20569 and n20823_not n20824_not ; f[83]
g20570 and n20569_not n20813_not ; n20826
g20571 and n20566_not n20826_not ; n20827
g20572 and b[63] n2048 ; n20828
g20573 and b[61] n2198 ; n20829
g20574 and b[62] n2043 ; n20830
g20575 and n20829_not n20830_not ; n20831
g20576 and n20828_not n20831 ; n20832
g20577 and n2051 n13771 ; n20833
g20578 and n20832 n20833_not ; n20834
g20579 and a[23] n20834_not ; n20835
g20580 and a[23] n20835_not ; n20836
g20581 and n20834_not n20835_not ; n20837
g20582 and n20836_not n20837_not ; n20838
g20583 and n20827_not n20838_not ; n20839
g20584 and n20827_not n20839_not ; n20840
g20585 and n20838_not n20839_not ; n20841
g20586 and n20840_not n20841_not ; n20842
g20587 and b[60] n2539 ; n20843
g20588 and b[58] n2685 ; n20844
g20589 and b[59] n2534 ; n20845
g20590 and n20844_not n20845_not ; n20846
g20591 and n20843_not n20846 ; n20847
g20592 and n2542 n12211 ; n20848
g20593 and n20847 n20848_not ; n20849
g20594 and a[26] n20849_not ; n20850
g20595 and a[26] n20850_not ; n20851
g20596 and n20849_not n20850_not ; n20852
g20597 and n20851_not n20852_not ; n20853
g20598 and n20583_not n20810_not ; n20854
g20599 and n20853 n20854 ; n20855
g20600 and n20853_not n20854_not ; n20856
g20601 and n20855_not n20856_not ; n20857
g20602 and n20600_not n20806_not ; n20858
g20603 and n20597_not n20858_not ; n20859
g20604 and b[57] n3050 ; n20860
g20605 and b[55] n3243 ; n20861
g20606 and b[56] n3045 ; n20862
g20607 and n20861_not n20862_not ; n20863
g20608 and n20860_not n20863 ; n20864
g20609 and n3053 n11410 ; n20865
g20610 and n20864 n20865_not ; n20866
g20611 and a[29] n20866_not ; n20867
g20612 and a[29] n20867_not ; n20868
g20613 and n20866_not n20867_not ; n20869
g20614 and n20868_not n20869_not ; n20870
g20615 and n20859_not n20870 ; n20871
g20616 and n20859 n20870_not ; n20872
g20617 and n20871_not n20872_not ; n20873
g20618 and b[54] n3638 ; n20874
g20619 and b[52] n3843 ; n20875
g20620 and b[53] n3633 ; n20876
g20621 and n20875_not n20876_not ; n20877
g20622 and n20874_not n20877 ; n20878
g20623 and n3641 n9998 ; n20879
g20624 and n20878 n20879_not ; n20880
g20625 and a[32] n20880_not ; n20881
g20626 and a[32] n20881_not ; n20882
g20627 and n20880_not n20881_not ; n20883
g20628 and n20882_not n20883_not ; n20884
g20629 and n20614_not n20802_not ; n20885
g20630 and n20884 n20885 ; n20886
g20631 and n20884_not n20885_not ; n20887
g20632 and n20886_not n20887_not ; n20888
g20633 and n20786_not n20799_not ; n20889
g20634 and n20742_not n20745_not ; n20890
g20635 and b[20] n13903 ; n20891
g20636 and b[21] n13488_not ; n20892
g20637 and n20891_not n20892_not ; n20893
g20638 and a[20]_not n20893_not ; n20894
g20639 and a[20] n20893 ; n20895
g20640 and n20894_not n20895_not ; n20896
g20641 and n20680_not n20896 ; n20897
g20642 and n20680 n20896_not ; n20898
g20643 and n20897_not n20898_not ; n20899
g20644 and b[24] n12668 ; n20900
g20645 and b[22] n13047 ; n20901
g20646 and b[23] n12663 ; n20902
g20647 and n20901_not n20902_not ; n20903
g20648 and n20900_not n20903 ; n20904
g20649 and n2458 n12671 ; n20905
g20650 and n20904 n20905_not ; n20906
g20651 and a[62] n20906_not ; n20907
g20652 and a[62] n20907_not ; n20908
g20653 and n20906_not n20907_not ; n20909
g20654 and n20908_not n20909_not ; n20910
g20655 and n20899 n20910_not ; n20911
g20656 and n20899 n20911_not ; n20912
g20657 and n20910_not n20911_not ; n20913
g20658 and n20912_not n20913_not ; n20914
g20659 and n20681_not n20695_not ; n20915
g20660 and n20914_not n20915_not ; n20916
g20661 and n20914_not n20916_not ; n20917
g20662 and n20915_not n20916_not ; n20918
g20663 and n20917_not n20918_not ; n20919
g20664 and b[27] n11531 ; n20920
g20665 and b[25] n11896 ; n20921
g20666 and b[26] n11526 ; n20922
g20667 and n20921_not n20922_not ; n20923
g20668 and n20920_not n20923 ; n20924
g20669 and n2990 n11534 ; n20925
g20670 and n20924 n20925_not ; n20926
g20671 and a[59] n20926_not ; n20927
g20672 and a[59] n20927_not ; n20928
g20673 and n20926_not n20927_not ; n20929
g20674 and n20928_not n20929_not ; n20930
g20675 and n20919_not n20930_not ; n20931
g20676 and n20919_not n20931_not ; n20932
g20677 and n20930_not n20931_not ; n20933
g20678 and n20932_not n20933_not ; n20934
g20679 and n20698_not n20701_not ; n20935
g20680 and n20934 n20935 ; n20936
g20681 and n20934_not n20935_not ; n20937
g20682 and n20936_not n20937_not ; n20938
g20683 and b[30] n10426 ; n20939
g20684 and b[28] n10796 ; n20940
g20685 and b[29] n10421 ; n20941
g20686 and n20940_not n20941_not ; n20942
g20687 and n20939_not n20942 ; n20943
g20688 and n3577 n10429 ; n20944
g20689 and n20943 n20944_not ; n20945
g20690 and a[56] n20945_not ; n20946
g20691 and a[56] n20946_not ; n20947
g20692 and n20945_not n20946_not ; n20948
g20693 and n20947_not n20948_not ; n20949
g20694 and n20938 n20949_not ; n20950
g20695 and n20938 n20950_not ; n20951
g20696 and n20949_not n20950_not ; n20952
g20697 and n20951_not n20952_not ; n20953
g20698 and n20704_not n20718_not ; n20954
g20699 and n20953 n20954 ; n20955
g20700 and n20953_not n20954_not ; n20956
g20701 and n20955_not n20956_not ; n20957
g20702 and b[33] n9339 ; n20958
g20703 and b[31] n9732 ; n20959
g20704 and b[32] n9334 ; n20960
g20705 and n20959_not n20960_not ; n20961
g20706 and n20958_not n20961 ; n20962
g20707 and n4223 n9342 ; n20963
g20708 and n20962 n20963_not ; n20964
g20709 and a[53] n20964_not ; n20965
g20710 and a[53] n20965_not ; n20966
g20711 and n20964_not n20965_not ; n20967
g20712 and n20966_not n20967_not ; n20968
g20713 and n20727_not n20738_not ; n20969
g20714 and n20724_not n20969_not ; n20970
g20715 and n20968_not n20970_not ; n20971
g20716 and n20968 n20970 ; n20972
g20717 and n20971_not n20972_not ; n20973
g20718 and n20957_not n20973 ; n20974
g20719 and n20957 n20973_not ; n20975
g20720 and n20974_not n20975_not ; n20976
g20721 and b[36] n8362 ; n20977
g20722 and b[34] n8715 ; n20978
g20723 and b[35] n8357 ; n20979
g20724 and n20978_not n20979_not ; n20980
g20725 and n20977_not n20980 ; n20981
g20726 and n4922 n8365 ; n20982
g20727 and n20981 n20982_not ; n20983
g20728 and a[50] n20983_not ; n20984
g20729 and a[50] n20984_not ; n20985
g20730 and n20983_not n20984_not ; n20986
g20731 and n20985_not n20986_not ; n20987
g20732 and n20976_not n20987_not ; n20988
g20733 and n20976 n20987 ; n20989
g20734 and n20988_not n20989_not ; n20990
g20735 and n20890 n20990_not ; n20991
g20736 and n20890_not n20990 ; n20992
g20737 and n20991_not n20992_not ; n20993
g20738 and b[39] n7446 ; n20994
g20739 and b[37] n7787 ; n20995
g20740 and b[38] n7441 ; n20996
g20741 and n20995_not n20996_not ; n20997
g20742 and n20994_not n20997 ; n20998
g20743 and n5451 n7449 ; n20999
g20744 and n20998 n20999_not ; n21000
g20745 and a[47] n21000_not ; n21001
g20746 and a[47] n21001_not ; n21002
g20747 and n21000_not n21001_not ; n21003
g20748 and n21002_not n21003_not ; n21004
g20749 and n20993 n21004_not ; n21005
g20750 and n20993 n21005_not ; n21006
g20751 and n21004_not n21005_not ; n21007
g20752 and n21006_not n21007_not ; n21008
g20753 and n20748_not n20751_not ; n21009
g20754 and n21008 n21009 ; n21010
g20755 and n21008_not n21009_not ; n21011
g20756 and n21010_not n21011_not ; n21012
g20757 and b[42] n6595 ; n21013
g20758 and b[40] n6902 ; n21014
g20759 and b[41] n6590 ; n21015
g20760 and n21014_not n21015_not ; n21016
g20761 and n21013_not n21016 ; n21017
g20762 and n6489 n6598 ; n21018
g20763 and n21017 n21018_not ; n21019
g20764 and a[44] n21019_not ; n21020
g20765 and a[44] n21020_not ; n21021
g20766 and n21019_not n21020_not ; n21022
g20767 and n21021_not n21022_not ; n21023
g20768 and n21012 n21023_not ; n21024
g20769 and n21012 n21024_not ; n21025
g20770 and n21023_not n21024_not ; n21026
g20771 and n21025_not n21026_not ; n21027
g20772 and n20754_not n20757_not ; n21028
g20773 and n21027 n21028 ; n21029
g20774 and n21027_not n21028_not ; n21030
g20775 and n21029_not n21030_not ; n21031
g20776 and b[45] n5777 ; n21032
g20777 and b[43] n6059 ; n21033
g20778 and b[44] n5772 ; n21034
g20779 and n21033_not n21034_not ; n21035
g20780 and n21032_not n21035 ; n21036
g20781 and n5780 n7361 ; n21037
g20782 and n21036 n21037_not ; n21038
g20783 and a[41] n21038_not ; n21039
g20784 and a[41] n21039_not ; n21040
g20785 and n21038_not n21039_not ; n21041
g20786 and n21040_not n21041_not ; n21042
g20787 and n21031 n21042_not ; n21043
g20788 and n21031 n21043_not ; n21044
g20789 and n21042_not n21043_not ; n21045
g20790 and n21044_not n21045_not ; n21046
g20791 and n20760_not n20763_not ; n21047
g20792 and n21046 n21047 ; n21048
g20793 and n21046_not n21047_not ; n21049
g20794 and n21048_not n21049_not ; n21050
g20795 and b[48] n5035 ; n21051
g20796 and b[46] n5277 ; n21052
g20797 and b[47] n5030 ; n21053
g20798 and n21052_not n21053_not ; n21054
g20799 and n21051_not n21054 ; n21055
g20800 and n5038 n8009 ; n21056
g20801 and n21055 n21056_not ; n21057
g20802 and a[38] n21057_not ; n21058
g20803 and a[38] n21058_not ; n21059
g20804 and n21057_not n21058_not ; n21060
g20805 and n21059_not n21060_not ; n21061
g20806 and n21050 n21061_not ; n21062
g20807 and n21050 n21062_not ; n21063
g20808 and n21061_not n21062_not ; n21064
g20809 and n21063_not n21064_not ; n21065
g20810 and n20766_not n20780_not ; n21066
g20811 and n21065 n21066 ; n21067
g20812 and n21065_not n21066_not ; n21068
g20813 and n21067_not n21068_not ; n21069
g20814 and b[51] n4287 ; n21070
g20815 and b[49] n4532 ; n21071
g20816 and b[50] n4282 ; n21072
g20817 and n21071_not n21072_not ; n21073
g20818 and n21070_not n21073 ; n21074
g20819 and n4290 n8976 ; n21075
g20820 and n21074 n21075_not ; n21076
g20821 and a[35] n21076_not ; n21077
g20822 and a[35] n21077_not ; n21078
g20823 and n21076_not n21077_not ; n21079
g20824 and n21078_not n21079_not ; n21080
g20825 and n21069 n21080_not ; n21081
g20826 and n21069_not n21080 ; n21082
g20827 and n20889_not n21082_not ; n21083
g20828 and n21081_not n21083 ; n21084
g20829 and n20889_not n21084_not ; n21085
g20830 and n21081_not n21084_not ; n21086
g20831 and n21082_not n21086 ; n21087
g20832 and n21085_not n21087_not ; n21088
g20833 and n20888 n21088_not ; n21089
g20834 and n20888_not n21088 ; n21090
g20835 and n20873_not n21090_not ; n21091
g20836 and n21089_not n21091 ; n21092
g20837 and n20873_not n21092_not ; n21093
g20838 and n21090_not n21092_not ; n21094
g20839 and n21089_not n21094 ; n21095
g20840 and n21093_not n21095_not ; n21096
g20841 and n20857 n21096_not ; n21097
g20842 and n20857_not n21096 ; n21098
g20843 and n20842_not n21098_not ; n21099
g20844 and n21097_not n21099 ; n21100
g20845 and n20842_not n21100_not ; n21101
g20846 and n21098_not n21100_not ; n21102
g20847 and n21097_not n21102 ; n21103
g20848 and n21101_not n21103_not ; n21104
g20849 and n20550_not n20817_not ; n21105
g20850 and n21104 n21105 ; n21106
g20851 and n21104_not n21105_not ; n21107
g20852 and n21106_not n21107_not ; n21108
g20853 and n20820_not n20823_not ; n21109
g20854 and n21108 n21109_not ; n21110
g20855 and n21108_not n21109 ; n21111
g20856 and n21110_not n21111_not ; f[84]
g20857 and n20856_not n21097_not ; n21113
g20858 and b[62] n2198 ; n21114
g20859 and b[63] n2043 ; n21115
g20860 and n21114_not n21115_not ; n21116
g20861 and n2051_not n21116 ; n21117
g20862 and n13800 n21116 ; n21118
g20863 and n21117_not n21118_not ; n21119
g20864 and a[23] n21119_not ; n21120
g20865 and a[23]_not n21119 ; n21121
g20866 and n21120_not n21121_not ; n21122
g20867 and n21113_not n21122_not ; n21123
g20868 and n21113 n21122 ; n21124
g20869 and n21123_not n21124_not ; n21125
g20870 and b[61] n2539 ; n21126
g20871 and b[59] n2685 ; n21127
g20872 and b[60] n2534 ; n21128
g20873 and n21127_not n21128_not ; n21129
g20874 and n21126_not n21129 ; n21130
g20875 and n2542 n12969 ; n21131
g20876 and n21130 n21131_not ; n21132
g20877 and a[26] n21132_not ; n21133
g20878 and a[26] n21133_not ; n21134
g20879 and n21132_not n21133_not ; n21135
g20880 and n21134_not n21135_not ; n21136
g20881 and n20859_not n20870_not ; n21137
g20882 and n21092_not n21137_not ; n21138
g20883 and n21136 n21138 ; n21139
g20884 and n21136_not n21138_not ; n21140
g20885 and n21139_not n21140_not ; n21141
g20886 and n20887_not n21089_not ; n21142
g20887 and b[58] n3050 ; n21143
g20888 and b[56] n3243 ; n21144
g20889 and b[57] n3045 ; n21145
g20890 and n21144_not n21145_not ; n21146
g20891 and n21143_not n21146 ; n21147
g20892 and n3053_not n21147 ; n21148
g20893 and n11436_not n21147 ; n21149
g20894 and n21148_not n21149_not ; n21150
g20895 and a[29] n21150_not ; n21151
g20896 and a[29]_not n21150 ; n21152
g20897 and n21151_not n21152_not ; n21153
g20898 and n21142_not n21153_not ; n21154
g20899 and n21142 n21153 ; n21155
g20900 and n21154_not n21155_not ; n21156
g20901 and b[55] n3638 ; n21157
g20902 and b[53] n3843 ; n21158
g20903 and b[54] n3633 ; n21159
g20904 and n21158_not n21159_not ; n21160
g20905 and n21157_not n21160 ; n21161
g20906 and n3641 n10684 ; n21162
g20907 and n21161 n21162_not ; n21163
g20908 and a[32] n21163_not ; n21164
g20909 and a[32] n21164_not ; n21165
g20910 and n21163_not n21164_not ; n21166
g20911 and n21165_not n21166_not ; n21167
g20912 and n21086_not n21167 ; n21168
g20913 and n21086 n21167_not ; n21169
g20914 and n21168_not n21169_not ; n21170
g20915 and b[43] n6595 ; n21171
g20916 and b[41] n6902 ; n21172
g20917 and b[42] n6590 ; n21173
g20918 and n21172_not n21173_not ; n21174
g20919 and n21171_not n21174 ; n21175
g20920 and n6515 n6598 ; n21176
g20921 and n21175 n21176_not ; n21177
g20922 and a[44] n21177_not ; n21178
g20923 and a[44] n21178_not ; n21179
g20924 and n21177_not n21178_not ; n21180
g20925 and n21179_not n21180_not ; n21181
g20926 and n21005_not n21011_not ; n21182
g20927 and b[40] n7446 ; n21183
g20928 and b[38] n7787 ; n21184
g20929 and b[39] n7441 ; n21185
g20930 and n21184_not n21185_not ; n21186
g20931 and n21183_not n21186 ; n21187
g20932 and n5955 n7449 ; n21188
g20933 and n21187 n21188_not ; n21189
g20934 and a[47] n21189_not ; n21190
g20935 and a[47] n21190_not ; n21191
g20936 and n21189_not n21190_not ; n21192
g20937 and n21191_not n21192_not ; n21193
g20938 and n20988_not n20992_not ; n21194
g20939 and n20931_not n20937_not ; n21195
g20940 and b[28] n11531 ; n21196
g20941 and b[26] n11896 ; n21197
g20942 and b[27] n11526 ; n21198
g20943 and n21197_not n21198_not ; n21199
g20944 and n21196_not n21199 ; n21200
g20945 and n3189 n11534 ; n21201
g20946 and n21200 n21201_not ; n21202
g20947 and a[59] n21202_not ; n21203
g20948 and a[59] n21203_not ; n21204
g20949 and n21202_not n21203_not ; n21205
g20950 and n21204_not n21205_not ; n21206
g20951 and n20911_not n20916_not ; n21207
g20952 and b[21] n13903 ; n21208
g20953 and b[22] n13488_not ; n21209
g20954 and n21208_not n21209_not ; n21210
g20955 and n20894_not n20897_not ; n21211
g20956 and n21210_not n21211 ; n21212
g20957 and n21210 n21211_not ; n21213
g20958 and n21212_not n21213_not ; n21214
g20959 and b[25] n12668 ; n21215
g20960 and b[23] n13047 ; n21216
g20961 and b[24] n12663 ; n21217
g20962 and n21216_not n21217_not ; n21218
g20963 and n21215_not n21218 ; n21219
g20964 and n12671_not n21219 ; n21220
g20965 and n2485_not n21219 ; n21221
g20966 and n21220_not n21221_not ; n21222
g20967 and a[62] n21222_not ; n21223
g20968 and a[62]_not n21222 ; n21224
g20969 and n21223_not n21224_not ; n21225
g20970 and n21214 n21225_not ; n21226
g20971 and n21214_not n21225 ; n21227
g20972 and n21226_not n21227_not ; n21228
g20973 and n21207_not n21228 ; n21229
g20974 and n21207 n21228_not ; n21230
g20975 and n21229_not n21230_not ; n21231
g20976 and n21206_not n21231 ; n21232
g20977 and n21206 n21231_not ; n21233
g20978 and n21232_not n21233_not ; n21234
g20979 and n21195_not n21234 ; n21235
g20980 and n21195 n21234_not ; n21236
g20981 and n21235_not n21236_not ; n21237
g20982 and b[31] n10426 ; n21238
g20983 and b[29] n10796 ; n21239
g20984 and b[30] n10421 ; n21240
g20985 and n21239_not n21240_not ; n21241
g20986 and n21238_not n21241 ; n21242
g20987 and n3796 n10429 ; n21243
g20988 and n21242 n21243_not ; n21244
g20989 and a[56] n21244_not ; n21245
g20990 and a[56] n21245_not ; n21246
g20991 and n21244_not n21245_not ; n21247
g20992 and n21246_not n21247_not ; n21248
g20993 and n21237 n21248_not ; n21249
g20994 and n21237 n21249_not ; n21250
g20995 and n21248_not n21249_not ; n21251
g20996 and n21250_not n21251_not ; n21252
g20997 and n20950_not n20956_not ; n21253
g20998 and n21252 n21253 ; n21254
g20999 and n21252_not n21253_not ; n21255
g21000 and n21254_not n21255_not ; n21256
g21001 and b[34] n9339 ; n21257
g21002 and b[32] n9732 ; n21258
g21003 and b[33] n9334 ; n21259
g21004 and n21258_not n21259_not ; n21260
g21005 and n21257_not n21260 ; n21261
g21006 and n4466 n9342 ; n21262
g21007 and n21261 n21262_not ; n21263
g21008 and a[53] n21263_not ; n21264
g21009 and a[53] n21264_not ; n21265
g21010 and n21263_not n21264_not ; n21266
g21011 and n21265_not n21266_not ; n21267
g21012 and n21256 n21267_not ; n21268
g21013 and n21256 n21268_not ; n21269
g21014 and n21267_not n21268_not ; n21270
g21015 and n21269_not n21270_not ; n21271
g21016 and n20957 n20973 ; n21272
g21017 and n20971_not n21272_not ; n21273
g21018 and n21271 n21273 ; n21274
g21019 and n21271_not n21273_not ; n21275
g21020 and n21274_not n21275_not ; n21276
g21021 and b[37] n8362 ; n21277
g21022 and b[35] n8715 ; n21278
g21023 and b[36] n8357 ; n21279
g21024 and n21278_not n21279_not ; n21280
g21025 and n21277_not n21280 ; n21281
g21026 and n5181 n8365 ; n21282
g21027 and n21281 n21282_not ; n21283
g21028 and a[50] n21283_not ; n21284
g21029 and a[50] n21284_not ; n21285
g21030 and n21283_not n21284_not ; n21286
g21031 and n21285_not n21286_not ; n21287
g21032 and n21276_not n21287 ; n21288
g21033 and n21276 n21287_not ; n21289
g21034 and n21288_not n21289_not ; n21290
g21035 and n21194_not n21290 ; n21291
g21036 and n21194_not n21291_not ; n21292
g21037 and n21290 n21291_not ; n21293
g21038 and n21292_not n21293_not ; n21294
g21039 and n21193_not n21294_not ; n21295
g21040 and n21193 n21293_not ; n21296
g21041 and n21292_not n21296 ; n21297
g21042 and n21295_not n21297_not ; n21298
g21043 and n21182_not n21298 ; n21299
g21044 and n21182 n21298_not ; n21300
g21045 and n21299_not n21300_not ; n21301
g21046 and n21181_not n21301 ; n21302
g21047 and n21301 n21302_not ; n21303
g21048 and n21181_not n21302_not ; n21304
g21049 and n21303_not n21304_not ; n21305
g21050 and n21024_not n21030_not ; n21306
g21051 and n21305 n21306 ; n21307
g21052 and n21305_not n21306_not ; n21308
g21053 and n21307_not n21308_not ; n21309
g21054 and b[46] n5777 ; n21310
g21055 and b[44] n6059 ; n21311
g21056 and b[45] n5772 ; n21312
g21057 and n21311_not n21312_not ; n21313
g21058 and n21310_not n21313 ; n21314
g21059 and n5780 n7677 ; n21315
g21060 and n21314 n21315_not ; n21316
g21061 and a[41] n21316_not ; n21317
g21062 and a[41] n21317_not ; n21318
g21063 and n21316_not n21317_not ; n21319
g21064 and n21318_not n21319_not ; n21320
g21065 and n21309 n21320_not ; n21321
g21066 and n21309 n21321_not ; n21322
g21067 and n21320_not n21321_not ; n21323
g21068 and n21322_not n21323_not ; n21324
g21069 and n21043_not n21049_not ; n21325
g21070 and n21324 n21325 ; n21326
g21071 and n21324_not n21325_not ; n21327
g21072 and n21326_not n21327_not ; n21328
g21073 and b[49] n5035 ; n21329
g21074 and b[47] n5277 ; n21330
g21075 and b[48] n5030 ; n21331
g21076 and n21330_not n21331_not ; n21332
g21077 and n21329_not n21332 ; n21333
g21078 and n5038 n8625 ; n21334
g21079 and n21333 n21334_not ; n21335
g21080 and a[38] n21335_not ; n21336
g21081 and a[38] n21336_not ; n21337
g21082 and n21335_not n21336_not ; n21338
g21083 and n21337_not n21338_not ; n21339
g21084 and n21328 n21339_not ; n21340
g21085 and n21328 n21340_not ; n21341
g21086 and n21339_not n21340_not ; n21342
g21087 and n21341_not n21342_not ; n21343
g21088 and n21062_not n21068_not ; n21344
g21089 and n21343 n21344 ; n21345
g21090 and n21343_not n21344_not ; n21346
g21091 and n21345_not n21346_not ; n21347
g21092 and b[52] n4287 ; n21348
g21093 and b[50] n4532 ; n21349
g21094 and b[51] n4282 ; n21350
g21095 and n21349_not n21350_not ; n21351
g21096 and n21348_not n21351 ; n21352
g21097 and n4290 n9628 ; n21353
g21098 and n21352 n21353_not ; n21354
g21099 and a[35] n21354_not ; n21355
g21100 and a[35] n21355_not ; n21356
g21101 and n21354_not n21355_not ; n21357
g21102 and n21356_not n21357_not ; n21358
g21103 and n21347 n21358_not ; n21359
g21104 and n21347 n21359_not ; n21360
g21105 and n21358_not n21359_not ; n21361
g21106 and n21360_not n21361_not ; n21362
g21107 and n21170_not n21362_not ; n21363
g21108 and n21170 n21362 ; n21364
g21109 and n21156 n21364_not ; n21365
g21110 and n21363_not n21365 ; n21366
g21111 and n21156 n21366_not ; n21367
g21112 and n21364_not n21366_not ; n21368
g21113 and n21363_not n21368 ; n21369
g21114 and n21367_not n21369_not ; n21370
g21115 and n21141 n21370_not ; n21371
g21116 and n21141_not n21370 ; n21372
g21117 and n21125 n21372_not ; n21373
g21118 and n21371_not n21373 ; n21374
g21119 and n21125 n21374_not ; n21375
g21120 and n21372_not n21374_not ; n21376
g21121 and n21371_not n21376 ; n21377
g21122 and n21375_not n21377_not ; n21378
g21123 and n20839_not n21100_not ; n21379
g21124 and n21378 n21379 ; n21380
g21125 and n21378_not n21379_not ; n21381
g21126 and n21380_not n21381_not ; n21382
g21127 and n21107_not n21110_not ; n21383
g21128 and n21382 n21383_not ; n21384
g21129 and n21382_not n21383 ; n21385
g21130 and n21384_not n21385_not ; f[85]
g21131 and n21381_not n21384_not ; n21387
g21132 and n21123_not n21374_not ; n21388
g21133 and n21140_not n21371_not ; n21389
g21134 and b[63] n2198 ; n21390
g21135 and n2051 n13797 ; n21391
g21136 and n21390_not n21391_not ; n21392
g21137 and a[23] n21392_not ; n21393
g21138 and a[23] n21393_not ; n21394
g21139 and n21392_not n21393_not ; n21395
g21140 and n21394_not n21395_not ; n21396
g21141 and n21389_not n21396_not ; n21397
g21142 and n21389_not n21397_not ; n21398
g21143 and n21396_not n21397_not ; n21399
g21144 and n21398_not n21399_not ; n21400
g21145 and b[62] n2539 ; n21401
g21146 and b[60] n2685 ; n21402
g21147 and b[61] n2534 ; n21403
g21148 and n21402_not n21403_not ; n21404
g21149 and n21401_not n21404 ; n21405
g21150 and n2542 n13370 ; n21406
g21151 and n21405 n21406_not ; n21407
g21152 and a[26] n21407_not ; n21408
g21153 and a[26] n21408_not ; n21409
g21154 and n21407_not n21408_not ; n21410
g21155 and n21409_not n21410_not ; n21411
g21156 and n21154_not n21366_not ; n21412
g21157 and n21411 n21412 ; n21413
g21158 and n21411_not n21412_not ; n21414
g21159 and n21413_not n21414_not ; n21415
g21160 and b[59] n3050 ; n21416
g21161 and b[57] n3243 ; n21417
g21162 and b[58] n3045 ; n21418
g21163 and n21417_not n21418_not ; n21419
g21164 and n21416_not n21419 ; n21420
g21165 and n3053 n12179 ; n21421
g21166 and n21420 n21421_not ; n21422
g21167 and a[29] n21422_not ; n21423
g21168 and a[29] n21423_not ; n21424
g21169 and n21422_not n21423_not ; n21425
g21170 and n21424_not n21425_not ; n21426
g21171 and n21086_not n21167_not ; n21427
g21172 and n21363_not n21427_not ; n21428
g21173 and n21426_not n21428_not ; n21429
g21174 and n21426_not n21429_not ; n21430
g21175 and n21428_not n21429_not ; n21431
g21176 and n21430_not n21431_not ; n21432
g21177 and b[56] n3638 ; n21433
g21178 and b[54] n3843 ; n21434
g21179 and b[55] n3633 ; n21435
g21180 and n21434_not n21435_not ; n21436
g21181 and n21433_not n21436 ; n21437
g21182 and n3641 n10708 ; n21438
g21183 and n21437 n21438_not ; n21439
g21184 and a[32] n21439_not ; n21440
g21185 and a[32] n21440_not ; n21441
g21186 and n21439_not n21440_not ; n21442
g21187 and n21441_not n21442_not ; n21443
g21188 and n21346_not n21359_not ; n21444
g21189 and n21443 n21444 ; n21445
g21190 and n21443_not n21444_not ; n21446
g21191 and n21445_not n21446_not ; n21447
g21192 and b[53] n4287 ; n21448
g21193 and b[51] n4532 ; n21449
g21194 and b[52] n4282 ; n21450
g21195 and n21449_not n21450_not ; n21451
g21196 and n21448_not n21451 ; n21452
g21197 and n4290 n9972 ; n21453
g21198 and n21452 n21453_not ; n21454
g21199 and a[35] n21454_not ; n21455
g21200 and a[35] n21455_not ; n21456
g21201 and n21454_not n21455_not ; n21457
g21202 and n21456_not n21457_not ; n21458
g21203 and n21327_not n21340_not ; n21459
g21204 and n21299_not n21302_not ; n21460
g21205 and b[44] n6595 ; n21461
g21206 and b[42] n6902 ; n21462
g21207 and b[43] n6590 ; n21463
g21208 and n21462_not n21463_not ; n21464
g21209 and n21461_not n21464 ; n21465
g21210 and n6598 n7072 ; n21466
g21211 and n21465 n21466_not ; n21467
g21212 and a[44] n21467_not ; n21468
g21213 and a[44] n21468_not ; n21469
g21214 and n21467_not n21468_not ; n21470
g21215 and n21469_not n21470_not ; n21471
g21216 and n21291_not n21295_not ; n21472
g21217 and n21255_not n21268_not ; n21473
g21218 and b[35] n9339 ; n21474
g21219 and b[33] n9732 ; n21475
g21220 and b[34] n9334 ; n21476
g21221 and n21475_not n21476_not ; n21477
g21222 and n21474_not n21477 ; n21478
g21223 and n4696 n9342 ; n21479
g21224 and n21478 n21479_not ; n21480
g21225 and a[53] n21480_not ; n21481
g21226 and a[53] n21481_not ; n21482
g21227 and n21480_not n21481_not ; n21483
g21228 and n21482_not n21483_not ; n21484
g21229 and n21235_not n21249_not ; n21485
g21230 and n21213_not n21226_not ; n21486
g21231 and b[22] n13903 ; n21487
g21232 and b[23] n13488_not ; n21488
g21233 and n21487_not n21488_not ; n21489
g21234 and n21210_not n21489 ; n21490
g21235 and n21210 n21489_not ; n21491
g21236 and n21490_not n21491_not ; n21492
g21237 and b[26] n12668 ; n21493
g21238 and b[24] n13047 ; n21494
g21239 and b[25] n12663 ; n21495
g21240 and n21494_not n21495_not ; n21496
g21241 and n21493_not n21496 ; n21497
g21242 and n12671_not n21497 ; n21498
g21243 and n2813_not n21497 ; n21499
g21244 and n21498_not n21499_not ; n21500
g21245 and a[62] n21500_not ; n21501
g21246 and a[62]_not n21500 ; n21502
g21247 and n21501_not n21502_not ; n21503
g21248 and n21492 n21503_not ; n21504
g21249 and n21492_not n21503 ; n21505
g21250 and n21504_not n21505_not ; n21506
g21251 and n21486_not n21506 ; n21507
g21252 and n21486 n21506_not ; n21508
g21253 and n21507_not n21508_not ; n21509
g21254 and b[29] n11531 ; n21510
g21255 and b[27] n11896 ; n21511
g21256 and b[28] n11526 ; n21512
g21257 and n21511_not n21512_not ; n21513
g21258 and n21510_not n21513 ; n21514
g21259 and n3383 n11534 ; n21515
g21260 and n21514 n21515_not ; n21516
g21261 and a[59] n21516_not ; n21517
g21262 and a[59] n21517_not ; n21518
g21263 and n21516_not n21517_not ; n21519
g21264 and n21518_not n21519_not ; n21520
g21265 and n21509 n21520_not ; n21521
g21266 and n21509 n21521_not ; n21522
g21267 and n21520_not n21521_not ; n21523
g21268 and n21522_not n21523_not ; n21524
g21269 and n21229_not n21232_not ; n21525
g21270 and n21524 n21525 ; n21526
g21271 and n21524_not n21525_not ; n21527
g21272 and n21526_not n21527_not ; n21528
g21273 and b[32] n10426 ; n21529
g21274 and b[30] n10796 ; n21530
g21275 and b[31] n10421 ; n21531
g21276 and n21530_not n21531_not ; n21532
g21277 and n21529_not n21532 ; n21533
g21278 and n4013 n10429 ; n21534
g21279 and n21533 n21534_not ; n21535
g21280 and a[56] n21535_not ; n21536
g21281 and a[56] n21536_not ; n21537
g21282 and n21535_not n21536_not ; n21538
g21283 and n21537_not n21538_not ; n21539
g21284 and n21528_not n21539 ; n21540
g21285 and n21528 n21539_not ; n21541
g21286 and n21540_not n21541_not ; n21542
g21287 and n21485_not n21542 ; n21543
g21288 and n21485 n21542_not ; n21544
g21289 and n21543_not n21544_not ; n21545
g21290 and n21484_not n21545 ; n21546
g21291 and n21484 n21545_not ; n21547
g21292 and n21546_not n21547_not ; n21548
g21293 and n21473_not n21548 ; n21549
g21294 and n21473 n21548_not ; n21550
g21295 and n21549_not n21550_not ; n21551
g21296 and b[38] n8362 ; n21552
g21297 and b[36] n8715 ; n21553
g21298 and b[37] n8357 ; n21554
g21299 and n21553_not n21554_not ; n21555
g21300 and n21552_not n21555 ; n21556
g21301 and n5205 n8365 ; n21557
g21302 and n21556 n21557_not ; n21558
g21303 and a[50] n21558_not ; n21559
g21304 and a[50] n21559_not ; n21560
g21305 and n21558_not n21559_not ; n21561
g21306 and n21560_not n21561_not ; n21562
g21307 and n21551 n21562_not ; n21563
g21308 and n21551 n21563_not ; n21564
g21309 and n21562_not n21563_not ; n21565
g21310 and n21564_not n21565_not ; n21566
g21311 and n21275_not n21289_not ; n21567
g21312 and n21566_not n21567_not ; n21568
g21313 and n21566_not n21568_not ; n21569
g21314 and n21567_not n21568_not ; n21570
g21315 and n21569_not n21570_not ; n21571
g21316 and b[41] n7446 ; n21572
g21317 and b[39] n7787 ; n21573
g21318 and b[40] n7441 ; n21574
g21319 and n21573_not n21574_not ; n21575
g21320 and n21572_not n21575 ; n21576
g21321 and n6219 n7449 ; n21577
g21322 and n21576 n21577_not ; n21578
g21323 and a[47] n21578_not ; n21579
g21324 and a[47] n21579_not ; n21580
g21325 and n21578_not n21579_not ; n21581
g21326 and n21580_not n21581_not ; n21582
g21327 and n21571_not n21582 ; n21583
g21328 and n21571 n21582_not ; n21584
g21329 and n21583_not n21584_not ; n21585
g21330 and n21472_not n21585_not ; n21586
g21331 and n21472 n21585 ; n21587
g21332 and n21586_not n21587_not ; n21588
g21333 and n21471_not n21588 ; n21589
g21334 and n21471 n21588_not ; n21590
g21335 and n21589_not n21590_not ; n21591
g21336 and n21460_not n21591 ; n21592
g21337 and n21460 n21591_not ; n21593
g21338 and n21592_not n21593_not ; n21594
g21339 and b[47] n5777 ; n21595
g21340 and b[45] n6059 ; n21596
g21341 and b[46] n5772 ; n21597
g21342 and n21596_not n21597_not ; n21598
g21343 and n21595_not n21598 ; n21599
g21344 and n5780 n7703 ; n21600
g21345 and n21599 n21600_not ; n21601
g21346 and a[41] n21601_not ; n21602
g21347 and a[41] n21602_not ; n21603
g21348 and n21601_not n21602_not ; n21604
g21349 and n21603_not n21604_not ; n21605
g21350 and n21594 n21605_not ; n21606
g21351 and n21594 n21606_not ; n21607
g21352 and n21605_not n21606_not ; n21608
g21353 and n21607_not n21608_not ; n21609
g21354 and n21308_not n21321_not ; n21610
g21355 and n21609 n21610 ; n21611
g21356 and n21609_not n21610_not ; n21612
g21357 and n21611_not n21612_not ; n21613
g21358 and b[50] n5035 ; n21614
g21359 and b[48] n5277 ; n21615
g21360 and b[49] n5030 ; n21616
g21361 and n21615_not n21616_not ; n21617
g21362 and n21614_not n21617 ; n21618
g21363 and n5038 n8949 ; n21619
g21364 and n21618 n21619_not ; n21620
g21365 and a[38] n21620_not ; n21621
g21366 and a[38] n21621_not ; n21622
g21367 and n21620_not n21621_not ; n21623
g21368 and n21622_not n21623_not ; n21624
g21369 and n21613_not n21624 ; n21625
g21370 and n21613 n21624_not ; n21626
g21371 and n21625_not n21626_not ; n21627
g21372 and n21459_not n21627 ; n21628
g21373 and n21459_not n21628_not ; n21629
g21374 and n21627 n21628_not ; n21630
g21375 and n21629_not n21630_not ; n21631
g21376 and n21458_not n21631_not ; n21632
g21377 and n21458_not n21632_not ; n21633
g21378 and n21631_not n21632_not ; n21634
g21379 and n21633_not n21634_not ; n21635
g21380 and n21447 n21635_not ; n21636
g21381 and n21447 n21636_not ; n21637
g21382 and n21635_not n21636_not ; n21638
g21383 and n21637_not n21638_not ; n21639
g21384 and n21432_not n21639 ; n21640
g21385 and n21432 n21639_not ; n21641
g21386 and n21640_not n21641_not ; n21642
g21387 and n21415 n21642_not ; n21643
g21388 and n21415 n21643_not ; n21644
g21389 and n21642_not n21643_not ; n21645
g21390 and n21644_not n21645_not ; n21646
g21391 and n21400_not n21646 ; n21647
g21392 and n21400 n21646_not ; n21648
g21393 and n21647_not n21648_not ; n21649
g21394 and n21388_not n21649_not ; n21650
g21395 and n21388_not n21650_not ; n21651
g21396 and n21649_not n21650_not ; n21652
g21397 and n21651_not n21652_not ; n21653
g21398 and n21387_not n21653_not ; n21654
g21399 and n21387 n21652_not ; n21655
g21400 and n21651_not n21655 ; n21656
g21401 and n21654_not n21656_not ; f[86]
g21402 and n21650_not n21654_not ; n21658
g21403 and n21400_not n21646_not ; n21659
g21404 and n21397_not n21659_not ; n21660
g21405 and n21414_not n21643_not ; n21661
g21406 and b[63] n2539 ; n21662
g21407 and b[61] n2685 ; n21663
g21408 and b[62] n2534 ; n21664
g21409 and n21663_not n21664_not ; n21665
g21410 and n21662_not n21665 ; n21666
g21411 and n2542 n13771 ; n21667
g21412 and n21666 n21667_not ; n21668
g21413 and a[26] n21668_not ; n21669
g21414 and a[26] n21669_not ; n21670
g21415 and n21668_not n21669_not ; n21671
g21416 and n21670_not n21671_not ; n21672
g21417 and n21661_not n21672_not ; n21673
g21418 and n21661_not n21673_not ; n21674
g21419 and n21672_not n21673_not ; n21675
g21420 and n21674_not n21675_not ; n21676
g21421 and n21432_not n21639_not ; n21677
g21422 and n21429_not n21677_not ; n21678
g21423 and b[60] n3050 ; n21679
g21424 and b[58] n3243 ; n21680
g21425 and b[59] n3045 ; n21681
g21426 and n21680_not n21681_not ; n21682
g21427 and n21679_not n21682 ; n21683
g21428 and n3053 n12211 ; n21684
g21429 and n21683 n21684_not ; n21685
g21430 and a[29] n21685_not ; n21686
g21431 and a[29] n21686_not ; n21687
g21432 and n21685_not n21686_not ; n21688
g21433 and n21687_not n21688_not ; n21689
g21434 and n21678_not n21689 ; n21690
g21435 and n21678 n21689_not ; n21691
g21436 and n21690_not n21691_not ; n21692
g21437 and b[57] n3638 ; n21693
g21438 and b[55] n3843 ; n21694
g21439 and b[56] n3633 ; n21695
g21440 and n21694_not n21695_not ; n21696
g21441 and n21693_not n21696 ; n21697
g21442 and n3641 n11410 ; n21698
g21443 and n21697 n21698_not ; n21699
g21444 and a[32] n21699_not ; n21700
g21445 and a[32] n21700_not ; n21701
g21446 and n21699_not n21700_not ; n21702
g21447 and n21701_not n21702_not ; n21703
g21448 and n21446_not n21636_not ; n21704
g21449 and n21703 n21704 ; n21705
g21450 and n21703_not n21704_not ; n21706
g21451 and n21705_not n21706_not ; n21707
g21452 and n21628_not n21632_not ; n21708
g21453 and n21612_not n21626_not ; n21709
g21454 and n21586_not n21589_not ; n21710
g21455 and n21571_not n21582_not ; n21711
g21456 and n21568_not n21711_not ; n21712
g21457 and b[36] n9339 ; n21713
g21458 and b[34] n9732 ; n21714
g21459 and b[35] n9334 ; n21715
g21460 and n21714_not n21715_not ; n21716
g21461 and n21713_not n21716 ; n21717
g21462 and n4922 n9342 ; n21718
g21463 and n21717 n21718_not ; n21719
g21464 and a[53] n21719_not ; n21720
g21465 and a[53] n21720_not ; n21721
g21466 and n21719_not n21720_not ; n21722
g21467 and n21721_not n21722_not ; n21723
g21468 and n21507_not n21521_not ; n21724
g21469 and n21490_not n21504_not ; n21725
g21470 and b[23] n13903 ; n21726
g21471 and b[24] n13488_not ; n21727
g21472 and n21726_not n21727_not ; n21728
g21473 and a[23]_not n21728_not ; n21729
g21474 and a[23] n21728 ; n21730
g21475 and n21729_not n21730_not ; n21731
g21476 and n21489_not n21731 ; n21732
g21477 and n21489 n21731_not ; n21733
g21478 and n21732_not n21733_not ; n21734
g21479 and b[27] n12668 ; n21735
g21480 and b[25] n13047 ; n21736
g21481 and b[26] n12663 ; n21737
g21482 and n21736_not n21737_not ; n21738
g21483 and n21735_not n21738 ; n21739
g21484 and n2990 n12671 ; n21740
g21485 and n21739 n21740_not ; n21741
g21486 and a[62] n21741_not ; n21742
g21487 and a[62] n21742_not ; n21743
g21488 and n21741_not n21742_not ; n21744
g21489 and n21743_not n21744_not ; n21745
g21490 and n21734 n21745_not ; n21746
g21491 and n21734 n21746_not ; n21747
g21492 and n21745_not n21746_not ; n21748
g21493 and n21747_not n21748_not ; n21749
g21494 and n21725_not n21749 ; n21750
g21495 and n21725 n21749_not ; n21751
g21496 and n21750_not n21751_not ; n21752
g21497 and b[30] n11531 ; n21753
g21498 and b[28] n11896 ; n21754
g21499 and b[29] n11526 ; n21755
g21500 and n21754_not n21755_not ; n21756
g21501 and n21753_not n21756 ; n21757
g21502 and n3577 n11534 ; n21758
g21503 and n21757 n21758_not ; n21759
g21504 and a[59] n21759_not ; n21760
g21505 and a[59] n21760_not ; n21761
g21506 and n21759_not n21760_not ; n21762
g21507 and n21761_not n21762_not ; n21763
g21508 and n21752_not n21763_not ; n21764
g21509 and n21752 n21763 ; n21765
g21510 and n21764_not n21765_not ; n21766
g21511 and n21724 n21766_not ; n21767
g21512 and n21724_not n21766 ; n21768
g21513 and n21767_not n21768_not ; n21769
g21514 and b[33] n10426 ; n21770
g21515 and b[31] n10796 ; n21771
g21516 and b[32] n10421 ; n21772
g21517 and n21771_not n21772_not ; n21773
g21518 and n21770_not n21773 ; n21774
g21519 and n4223 n10429 ; n21775
g21520 and n21774 n21775_not ; n21776
g21521 and a[56] n21776_not ; n21777
g21522 and a[56] n21777_not ; n21778
g21523 and n21776_not n21777_not ; n21779
g21524 and n21778_not n21779_not ; n21780
g21525 and n21527_not n21541_not ; n21781
g21526 and n21780_not n21781_not ; n21782
g21527 and n21780 n21781 ; n21783
g21528 and n21782_not n21783_not ; n21784
g21529 and n21769 n21784 ; n21785
g21530 and n21769_not n21784_not ; n21786
g21531 and n21785_not n21786_not ; n21787
g21532 and n21723_not n21787 ; n21788
g21533 and n21787 n21788_not ; n21789
g21534 and n21723_not n21788_not ; n21790
g21535 and n21789_not n21790_not ; n21791
g21536 and n21543_not n21546_not ; n21792
g21537 and n21791 n21792 ; n21793
g21538 and n21791_not n21792_not ; n21794
g21539 and n21793_not n21794_not ; n21795
g21540 and b[39] n8362 ; n21796
g21541 and b[37] n8715 ; n21797
g21542 and b[38] n8357 ; n21798
g21543 and n21797_not n21798_not ; n21799
g21544 and n21796_not n21799 ; n21800
g21545 and n5451 n8365 ; n21801
g21546 and n21800 n21801_not ; n21802
g21547 and a[50] n21802_not ; n21803
g21548 and a[50] n21803_not ; n21804
g21549 and n21802_not n21803_not ; n21805
g21550 and n21804_not n21805_not ; n21806
g21551 and n21795 n21806_not ; n21807
g21552 and n21795 n21807_not ; n21808
g21553 and n21806_not n21807_not ; n21809
g21554 and n21808_not n21809_not ; n21810
g21555 and n21549_not n21563_not ; n21811
g21556 and n21810 n21811 ; n21812
g21557 and n21810_not n21811_not ; n21813
g21558 and n21812_not n21813_not ; n21814
g21559 and b[42] n7446 ; n21815
g21560 and b[40] n7787 ; n21816
g21561 and b[41] n7441 ; n21817
g21562 and n21816_not n21817_not ; n21818
g21563 and n21815_not n21818 ; n21819
g21564 and n6489 n7449 ; n21820
g21565 and n21819 n21820_not ; n21821
g21566 and a[47] n21821_not ; n21822
g21567 and a[47] n21822_not ; n21823
g21568 and n21821_not n21822_not ; n21824
g21569 and n21823_not n21824_not ; n21825
g21570 and n21814 n21825_not ; n21826
g21571 and n21814 n21826_not ; n21827
g21572 and n21825_not n21826_not ; n21828
g21573 and n21827_not n21828_not ; n21829
g21574 and n21712_not n21829 ; n21830
g21575 and n21712 n21829_not ; n21831
g21576 and n21830_not n21831_not ; n21832
g21577 and b[45] n6595 ; n21833
g21578 and b[43] n6902 ; n21834
g21579 and b[44] n6590 ; n21835
g21580 and n21834_not n21835_not ; n21836
g21581 and n21833_not n21836 ; n21837
g21582 and n6598 n7361 ; n21838
g21583 and n21837 n21838_not ; n21839
g21584 and a[44] n21839_not ; n21840
g21585 and a[44] n21840_not ; n21841
g21586 and n21839_not n21840_not ; n21842
g21587 and n21841_not n21842_not ; n21843
g21588 and n21832_not n21843_not ; n21844
g21589 and n21832 n21843 ; n21845
g21590 and n21844_not n21845_not ; n21846
g21591 and n21710 n21846_not ; n21847
g21592 and n21710_not n21846 ; n21848
g21593 and n21847_not n21848_not ; n21849
g21594 and b[48] n5777 ; n21850
g21595 and b[46] n6059 ; n21851
g21596 and b[47] n5772 ; n21852
g21597 and n21851_not n21852_not ; n21853
g21598 and n21850_not n21853 ; n21854
g21599 and n5780 n8009 ; n21855
g21600 and n21854 n21855_not ; n21856
g21601 and a[41] n21856_not ; n21857
g21602 and a[41] n21857_not ; n21858
g21603 and n21856_not n21857_not ; n21859
g21604 and n21858_not n21859_not ; n21860
g21605 and n21849 n21860_not ; n21861
g21606 and n21849 n21861_not ; n21862
g21607 and n21860_not n21861_not ; n21863
g21608 and n21862_not n21863_not ; n21864
g21609 and n21592_not n21606_not ; n21865
g21610 and n21864 n21865 ; n21866
g21611 and n21864_not n21865_not ; n21867
g21612 and n21866_not n21867_not ; n21868
g21613 and b[51] n5035 ; n21869
g21614 and b[49] n5277 ; n21870
g21615 and b[50] n5030 ; n21871
g21616 and n21870_not n21871_not ; n21872
g21617 and n21869_not n21872 ; n21873
g21618 and n5038 n8976 ; n21874
g21619 and n21873 n21874_not ; n21875
g21620 and a[38] n21875_not ; n21876
g21621 and a[38] n21876_not ; n21877
g21622 and n21875_not n21876_not ; n21878
g21623 and n21877_not n21878_not ; n21879
g21624 and n21868 n21879_not ; n21880
g21625 and n21868_not n21879 ; n21881
g21626 and n21709_not n21881_not ; n21882
g21627 and n21880_not n21882 ; n21883
g21628 and n21709_not n21883_not ; n21884
g21629 and n21880_not n21883_not ; n21885
g21630 and n21881_not n21885 ; n21886
g21631 and n21884_not n21886_not ; n21887
g21632 and b[54] n4287 ; n21888
g21633 and b[52] n4532 ; n21889
g21634 and b[53] n4282 ; n21890
g21635 and n21889_not n21890_not ; n21891
g21636 and n21888_not n21891 ; n21892
g21637 and n4290 n9998 ; n21893
g21638 and n21892 n21893_not ; n21894
g21639 and a[35] n21894_not ; n21895
g21640 and a[35] n21895_not ; n21896
g21641 and n21894_not n21895_not ; n21897
g21642 and n21896_not n21897_not ; n21898
g21643 and n21887 n21898 ; n21899
g21644 and n21887_not n21898_not ; n21900
g21645 and n21899_not n21900_not ; n21901
g21646 and n21708_not n21901 ; n21902
g21647 and n21708 n21901_not ; n21903
g21648 and n21902_not n21903_not ; n21904
g21649 and n21707 n21904 ; n21905
g21650 and n21707_not n21904_not ; n21906
g21651 and n21692_not n21906_not ; n21907
g21652 and n21905_not n21907 ; n21908
g21653 and n21692_not n21908_not ; n21909
g21654 and n21906_not n21908_not ; n21910
g21655 and n21905_not n21910 ; n21911
g21656 and n21909_not n21911_not ; n21912
g21657 and n21676_not n21912 ; n21913
g21658 and n21676 n21912_not ; n21914
g21659 and n21913_not n21914_not ; n21915
g21660 and n21660_not n21915_not ; n21916
g21661 and n21660_not n21916_not ; n21917
g21662 and n21915_not n21916_not ; n21918
g21663 and n21917_not n21918_not ; n21919
g21664 and n21658_not n21919_not ; n21920
g21665 and n21658 n21918_not ; n21921
g21666 and n21917_not n21921 ; n21922
g21667 and n21920_not n21922_not ; f[87]
g21668 and n21916_not n21920_not ; n21924
g21669 and n21676_not n21912_not ; n21925
g21670 and n21673_not n21925_not ; n21926
g21671 and b[61] n3050 ; n21927
g21672 and b[59] n3243 ; n21928
g21673 and b[60] n3045 ; n21929
g21674 and n21928_not n21929_not ; n21930
g21675 and n21927_not n21930 ; n21931
g21676 and n3053 n12969 ; n21932
g21677 and n21931 n21932_not ; n21933
g21678 and a[29] n21933_not ; n21934
g21679 and a[29] n21934_not ; n21935
g21680 and n21933_not n21934_not ; n21936
g21681 and n21935_not n21936_not ; n21937
g21682 and n21706_not n21905_not ; n21938
g21683 and n21937_not n21938_not ; n21939
g21684 and n21937_not n21939_not ; n21940
g21685 and n21938_not n21939_not ; n21941
g21686 and n21940_not n21941_not ; n21942
g21687 and n21900_not n21902_not ; n21943
g21688 and b[58] n3638 ; n21944
g21689 and b[56] n3843 ; n21945
g21690 and b[57] n3633 ; n21946
g21691 and n21945_not n21946_not ; n21947
g21692 and n21944_not n21947 ; n21948
g21693 and n3641_not n21948 ; n21949
g21694 and n11436_not n21948 ; n21950
g21695 and n21949_not n21950_not ; n21951
g21696 and a[32] n21951_not ; n21952
g21697 and a[32]_not n21951 ; n21953
g21698 and n21952_not n21953_not ; n21954
g21699 and n21943_not n21954_not ; n21955
g21700 and n21943 n21954 ; n21956
g21701 and n21955_not n21956_not ; n21957
g21702 and b[43] n7446 ; n21958
g21703 and b[41] n7787 ; n21959
g21704 and b[42] n7441 ; n21960
g21705 and n21959_not n21960_not ; n21961
g21706 and n21958_not n21961 ; n21962
g21707 and n6515 n7449 ; n21963
g21708 and n21962 n21963_not ; n21964
g21709 and a[47] n21964_not ; n21965
g21710 and a[47] n21965_not ; n21966
g21711 and n21964_not n21965_not ; n21967
g21712 and n21966_not n21967_not ; n21968
g21713 and n21807_not n21813_not ; n21969
g21714 and b[40] n8362 ; n21970
g21715 and b[38] n8715 ; n21971
g21716 and b[39] n8357 ; n21972
g21717 and n21971_not n21972_not ; n21973
g21718 and n21970_not n21973 ; n21974
g21719 and n5955 n8365 ; n21975
g21720 and n21974 n21975_not ; n21976
g21721 and a[50] n21976_not ; n21977
g21722 and a[50] n21977_not ; n21978
g21723 and n21976_not n21977_not ; n21979
g21724 and n21978_not n21979_not ; n21980
g21725 and n21788_not n21794_not ; n21981
g21726 and n21725_not n21749_not ; n21982
g21727 and n21746_not n21982_not ; n21983
g21728 and b[24] n13903 ; n21984
g21729 and b[25] n13488_not ; n21985
g21730 and n21984_not n21985_not ; n21986
g21731 and n21729_not n21732_not ; n21987
g21732 and n21986_not n21987 ; n21988
g21733 and n21986 n21987_not ; n21989
g21734 and n21988_not n21989_not ; n21990
g21735 and b[28] n12668 ; n21991
g21736 and b[26] n13047 ; n21992
g21737 and b[27] n12663 ; n21993
g21738 and n21992_not n21993_not ; n21994
g21739 and n21991_not n21994 ; n21995
g21740 and n12671_not n21995 ; n21996
g21741 and n3189_not n21995 ; n21997
g21742 and n21996_not n21997_not ; n21998
g21743 and a[62] n21998_not ; n21999
g21744 and a[62]_not n21998 ; n22000
g21745 and n21999_not n22000_not ; n22001
g21746 and n21990 n22001_not ; n22002
g21747 and n21990_not n22001 ; n22003
g21748 and n22002_not n22003_not ; n22004
g21749 and n21983_not n22004 ; n22005
g21750 and n21983 n22004_not ; n22006
g21751 and n22005_not n22006_not ; n22007
g21752 and b[31] n11531 ; n22008
g21753 and b[29] n11896 ; n22009
g21754 and b[30] n11526 ; n22010
g21755 and n22009_not n22010_not ; n22011
g21756 and n22008_not n22011 ; n22012
g21757 and n3796 n11534 ; n22013
g21758 and n22012 n22013_not ; n22014
g21759 and a[59] n22014_not ; n22015
g21760 and a[59] n22015_not ; n22016
g21761 and n22014_not n22015_not ; n22017
g21762 and n22016_not n22017_not ; n22018
g21763 and n22007 n22018_not ; n22019
g21764 and n22007 n22019_not ; n22020
g21765 and n22018_not n22019_not ; n22021
g21766 and n22020_not n22021_not ; n22022
g21767 and n21764_not n21768_not ; n22023
g21768 and n22022 n22023 ; n22024
g21769 and n22022_not n22023_not ; n22025
g21770 and n22024_not n22025_not ; n22026
g21771 and b[34] n10426 ; n22027
g21772 and b[32] n10796 ; n22028
g21773 and b[33] n10421 ; n22029
g21774 and n22028_not n22029_not ; n22030
g21775 and n22027_not n22030 ; n22031
g21776 and n4466 n10429 ; n22032
g21777 and n22031 n22032_not ; n22033
g21778 and a[56] n22033_not ; n22034
g21779 and a[56] n22034_not ; n22035
g21780 and n22033_not n22034_not ; n22036
g21781 and n22035_not n22036_not ; n22037
g21782 and n22026 n22037_not ; n22038
g21783 and n22026 n22038_not ; n22039
g21784 and n22037_not n22038_not ; n22040
g21785 and n22039_not n22040_not ; n22041
g21786 and n21782_not n21785_not ; n22042
g21787 and n22041 n22042 ; n22043
g21788 and n22041_not n22042_not ; n22044
g21789 and n22043_not n22044_not ; n22045
g21790 and b[37] n9339 ; n22046
g21791 and b[35] n9732 ; n22047
g21792 and b[36] n9334 ; n22048
g21793 and n22047_not n22048_not ; n22049
g21794 and n22046_not n22049 ; n22050
g21795 and n5181 n9342 ; n22051
g21796 and n22050 n22051_not ; n22052
g21797 and a[53] n22052_not ; n22053
g21798 and a[53] n22053_not ; n22054
g21799 and n22052_not n22053_not ; n22055
g21800 and n22054_not n22055_not ; n22056
g21801 and n22045_not n22056 ; n22057
g21802 and n22045 n22056_not ; n22058
g21803 and n22057_not n22058_not ; n22059
g21804 and n21981_not n22059 ; n22060
g21805 and n21981_not n22060_not ; n22061
g21806 and n22059 n22060_not ; n22062
g21807 and n22061_not n22062_not ; n22063
g21808 and n21980_not n22063_not ; n22064
g21809 and n21980 n22062_not ; n22065
g21810 and n22061_not n22065 ; n22066
g21811 and n22064_not n22066_not ; n22067
g21812 and n21969_not n22067 ; n22068
g21813 and n21969 n22067_not ; n22069
g21814 and n22068_not n22069_not ; n22070
g21815 and n21968_not n22070 ; n22071
g21816 and n22070 n22071_not ; n22072
g21817 and n21968_not n22071_not ; n22073
g21818 and n22072_not n22073_not ; n22074
g21819 and n21712_not n21829_not ; n22075
g21820 and n21826_not n22075_not ; n22076
g21821 and n22074 n22076 ; n22077
g21822 and n22074_not n22076_not ; n22078
g21823 and n22077_not n22078_not ; n22079
g21824 and b[46] n6595 ; n22080
g21825 and b[44] n6902 ; n22081
g21826 and b[45] n6590 ; n22082
g21827 and n22081_not n22082_not ; n22083
g21828 and n22080_not n22083 ; n22084
g21829 and n6598 n7677 ; n22085
g21830 and n22084 n22085_not ; n22086
g21831 and a[44] n22086_not ; n22087
g21832 and a[44] n22087_not ; n22088
g21833 and n22086_not n22087_not ; n22089
g21834 and n22088_not n22089_not ; n22090
g21835 and n22079 n22090_not ; n22091
g21836 and n22079 n22091_not ; n22092
g21837 and n22090_not n22091_not ; n22093
g21838 and n22092_not n22093_not ; n22094
g21839 and n21844_not n21848_not ; n22095
g21840 and n22094 n22095 ; n22096
g21841 and n22094_not n22095_not ; n22097
g21842 and n22096_not n22097_not ; n22098
g21843 and b[49] n5777 ; n22099
g21844 and b[47] n6059 ; n22100
g21845 and b[48] n5772 ; n22101
g21846 and n22100_not n22101_not ; n22102
g21847 and n22099_not n22102 ; n22103
g21848 and n5780 n8625 ; n22104
g21849 and n22103 n22104_not ; n22105
g21850 and a[41] n22105_not ; n22106
g21851 and a[41] n22106_not ; n22107
g21852 and n22105_not n22106_not ; n22108
g21853 and n22107_not n22108_not ; n22109
g21854 and n22098 n22109_not ; n22110
g21855 and n22098 n22110_not ; n22111
g21856 and n22109_not n22110_not ; n22112
g21857 and n22111_not n22112_not ; n22113
g21858 and n21861_not n21867_not ; n22114
g21859 and n22113 n22114 ; n22115
g21860 and n22113_not n22114_not ; n22116
g21861 and n22115_not n22116_not ; n22117
g21862 and b[52] n5035 ; n22118
g21863 and b[50] n5277 ; n22119
g21864 and b[51] n5030 ; n22120
g21865 and n22119_not n22120_not ; n22121
g21866 and n22118_not n22121 ; n22122
g21867 and n5038 n9628 ; n22123
g21868 and n22122 n22123_not ; n22124
g21869 and a[38] n22124_not ; n22125
g21870 and a[38] n22125_not ; n22126
g21871 and n22124_not n22125_not ; n22127
g21872 and n22126_not n22127_not ; n22128
g21873 and n22117 n22128_not ; n22129
g21874 and n22117 n22129_not ; n22130
g21875 and n22128_not n22129_not ; n22131
g21876 and n22130_not n22131_not ; n22132
g21877 and n21885_not n22132 ; n22133
g21878 and n21885 n22132_not ; n22134
g21879 and n22133_not n22134_not ; n22135
g21880 and b[55] n4287 ; n22136
g21881 and b[53] n4532 ; n22137
g21882 and b[54] n4282 ; n22138
g21883 and n22137_not n22138_not ; n22139
g21884 and n22136_not n22139 ; n22140
g21885 and n4290 n10684 ; n22141
g21886 and n22140 n22141_not ; n22142
g21887 and a[35] n22142_not ; n22143
g21888 and a[35] n22143_not ; n22144
g21889 and n22142_not n22143_not ; n22145
g21890 and n22144_not n22145_not ; n22146
g21891 and n22135_not n22146_not ; n22147
g21892 and n22135 n22146 ; n22148
g21893 and n22147_not n22148_not ; n22149
g21894 and n21957 n22149 ; n22150
g21895 and n21957_not n22149_not ; n22151
g21896 and n22150_not n22151_not ; n22152
g21897 and n21942_not n22152 ; n22153
g21898 and n21942_not n22153_not ; n22154
g21899 and n22152 n22153_not ; n22155
g21900 and n22154_not n22155_not ; n22156
g21901 and n21678_not n21689_not ; n22157
g21902 and n21908_not n22157_not ; n22158
g21903 and b[62] n2685 ; n22159
g21904 and b[63] n2534 ; n22160
g21905 and n22159_not n22160_not ; n22161
g21906 and n2542_not n22161 ; n22162
g21907 and n13800 n22161 ; n22163
g21908 and n22162_not n22163_not ; n22164
g21909 and a[26] n22164_not ; n22165
g21910 and a[26]_not n22164 ; n22166
g21911 and n22165_not n22166_not ; n22167
g21912 and n22158_not n22167_not ; n22168
g21913 and n22158_not n22168_not ; n22169
g21914 and n22167_not n22168_not ; n22170
g21915 and n22169_not n22170_not ; n22171
g21916 and n22156_not n22171_not ; n22172
g21917 and n22156 n22170_not ; n22173
g21918 and n22169_not n22173 ; n22174
g21919 and n22172_not n22174_not ; n22175
g21920 and n21926_not n22175 ; n22176
g21921 and n21926_not n22176_not ; n22177
g21922 and n22175 n22176_not ; n22178
g21923 and n22177_not n22178_not ; n22179
g21924 and n21924_not n22179_not ; n22180
g21925 and n21924 n22178_not ; n22181
g21926 and n22177_not n22181 ; n22182
g21927 and n22180_not n22182_not ; f[88]
g21928 and n22176_not n22180_not ; n22184
g21929 and n22168_not n22172_not ; n22185
g21930 and n21939_not n22153_not ; n22186
g21931 and b[63] n2685 ; n22187
g21932 and n2542 n13797 ; n22188
g21933 and n22187_not n22188_not ; n22189
g21934 and a[26] n22189_not ; n22190
g21935 and a[26] n22190_not ; n22191
g21936 and n22189_not n22190_not ; n22192
g21937 and n22191_not n22192_not ; n22193
g21938 and n22186_not n22193_not ; n22194
g21939 and n22186_not n22194_not ; n22195
g21940 and n22193_not n22194_not ; n22196
g21941 and n22195_not n22196_not ; n22197
g21942 and b[62] n3050 ; n22198
g21943 and b[60] n3243 ; n22199
g21944 and b[61] n3045 ; n22200
g21945 and n22199_not n22200_not ; n22201
g21946 and n22198_not n22201 ; n22202
g21947 and n3053 n13370 ; n22203
g21948 and n22202 n22203_not ; n22204
g21949 and a[29] n22204_not ; n22205
g21950 and a[29] n22205_not ; n22206
g21951 and n22204_not n22205_not ; n22207
g21952 and n22206_not n22207_not ; n22208
g21953 and n21955_not n22150_not ; n22209
g21954 and n22208 n22209 ; n22210
g21955 and n22208_not n22209_not ; n22211
g21956 and n22210_not n22211_not ; n22212
g21957 and b[59] n3638 ; n22213
g21958 and b[57] n3843 ; n22214
g21959 and b[58] n3633 ; n22215
g21960 and n22214_not n22215_not ; n22216
g21961 and n22213_not n22216 ; n22217
g21962 and n3641 n12179 ; n22218
g21963 and n22217 n22218_not ; n22219
g21964 and a[32] n22219_not ; n22220
g21965 and a[32] n22220_not ; n22221
g21966 and n22219_not n22220_not ; n22222
g21967 and n22221_not n22222_not ; n22223
g21968 and n21885_not n22132_not ; n22224
g21969 and n22147_not n22224_not ; n22225
g21970 and n22223 n22225 ; n22226
g21971 and n22223_not n22225_not ; n22227
g21972 and n22226_not n22227_not ; n22228
g21973 and b[56] n4287 ; n22229
g21974 and b[54] n4532 ; n22230
g21975 and b[55] n4282 ; n22231
g21976 and n22230_not n22231_not ; n22232
g21977 and n22229_not n22232 ; n22233
g21978 and n4290 n10708 ; n22234
g21979 and n22233 n22234_not ; n22235
g21980 and a[35] n22235_not ; n22236
g21981 and a[35] n22236_not ; n22237
g21982 and n22235_not n22236_not ; n22238
g21983 and n22237_not n22238_not ; n22239
g21984 and n22116_not n22129_not ; n22240
g21985 and b[53] n5035 ; n22241
g21986 and b[51] n5277 ; n22242
g21987 and b[52] n5030 ; n22243
g21988 and n22242_not n22243_not ; n22244
g21989 and n22241_not n22244 ; n22245
g21990 and n5038 n9972 ; n22246
g21991 and n22245 n22246_not ; n22247
g21992 and a[38] n22247_not ; n22248
g21993 and a[38] n22248_not ; n22249
g21994 and n22247_not n22248_not ; n22250
g21995 and n22249_not n22250_not ; n22251
g21996 and n22097_not n22110_not ; n22252
g21997 and n22068_not n22071_not ; n22253
g21998 and b[44] n7446 ; n22254
g21999 and b[42] n7787 ; n22255
g22000 and b[43] n7441 ; n22256
g22001 and n22255_not n22256_not ; n22257
g22002 and n22254_not n22257 ; n22258
g22003 and n7072 n7449 ; n22259
g22004 and n22258 n22259_not ; n22260
g22005 and a[47] n22260_not ; n22261
g22006 and a[47] n22261_not ; n22262
g22007 and n22260_not n22261_not ; n22263
g22008 and n22262_not n22263_not ; n22264
g22009 and n22060_not n22064_not ; n22265
g22010 and n22025_not n22038_not ; n22266
g22011 and b[35] n10426 ; n22267
g22012 and b[33] n10796 ; n22268
g22013 and b[34] n10421 ; n22269
g22014 and n22268_not n22269_not ; n22270
g22015 and n22267_not n22270 ; n22271
g22016 and n4696 n10429 ; n22272
g22017 and n22271 n22272_not ; n22273
g22018 and a[56] n22273_not ; n22274
g22019 and a[56] n22274_not ; n22275
g22020 and n22273_not n22274_not ; n22276
g22021 and n22275_not n22276_not ; n22277
g22022 and n22005_not n22019_not ; n22278
g22023 and b[32] n11531 ; n22279
g22024 and b[30] n11896 ; n22280
g22025 and b[31] n11526 ; n22281
g22026 and n22280_not n22281_not ; n22282
g22027 and n22279_not n22282 ; n22283
g22028 and n4013 n11534 ; n22284
g22029 and n22283 n22284_not ; n22285
g22030 and a[59] n22285_not ; n22286
g22031 and a[59] n22286_not ; n22287
g22032 and n22285_not n22286_not ; n22288
g22033 and n22287_not n22288_not ; n22289
g22034 and n21989_not n22002_not ; n22290
g22035 and b[25] n13903 ; n22291
g22036 and b[26] n13488_not ; n22292
g22037 and n22291_not n22292_not ; n22293
g22038 and n21986_not n22293 ; n22294
g22039 and n21986 n22293_not ; n22295
g22040 and n22294_not n22295_not ; n22296
g22041 and b[29] n12668 ; n22297
g22042 and b[27] n13047 ; n22298
g22043 and b[28] n12663 ; n22299
g22044 and n22298_not n22299_not ; n22300
g22045 and n22297_not n22300 ; n22301
g22046 and n12671_not n22301 ; n22302
g22047 and n3383_not n22301 ; n22303
g22048 and n22302_not n22303_not ; n22304
g22049 and a[62] n22304_not ; n22305
g22050 and a[62]_not n22304 ; n22306
g22051 and n22305_not n22306_not ; n22307
g22052 and n22296 n22307_not ; n22308
g22053 and n22296_not n22307 ; n22309
g22054 and n22308_not n22309_not ; n22310
g22055 and n22290_not n22310 ; n22311
g22056 and n22290 n22310_not ; n22312
g22057 and n22311_not n22312_not ; n22313
g22058 and n22289_not n22313 ; n22314
g22059 and n22289 n22313_not ; n22315
g22060 and n22314_not n22315_not ; n22316
g22061 and n22278_not n22316 ; n22317
g22062 and n22278 n22316_not ; n22318
g22063 and n22317_not n22318_not ; n22319
g22064 and n22277_not n22319 ; n22320
g22065 and n22277 n22319_not ; n22321
g22066 and n22320_not n22321_not ; n22322
g22067 and n22266_not n22322 ; n22323
g22068 and n22266 n22322_not ; n22324
g22069 and n22323_not n22324_not ; n22325
g22070 and b[38] n9339 ; n22326
g22071 and b[36] n9732 ; n22327
g22072 and b[37] n9334 ; n22328
g22073 and n22327_not n22328_not ; n22329
g22074 and n22326_not n22329 ; n22330
g22075 and n5205 n9342 ; n22331
g22076 and n22330 n22331_not ; n22332
g22077 and a[53] n22332_not ; n22333
g22078 and a[53] n22333_not ; n22334
g22079 and n22332_not n22333_not ; n22335
g22080 and n22334_not n22335_not ; n22336
g22081 and n22325 n22336_not ; n22337
g22082 and n22325 n22337_not ; n22338
g22083 and n22336_not n22337_not ; n22339
g22084 and n22338_not n22339_not ; n22340
g22085 and n22044_not n22058_not ; n22341
g22086 and n22340_not n22341_not ; n22342
g22087 and n22340_not n22342_not ; n22343
g22088 and n22341_not n22342_not ; n22344
g22089 and n22343_not n22344_not ; n22345
g22090 and b[41] n8362 ; n22346
g22091 and b[39] n8715 ; n22347
g22092 and b[40] n8357 ; n22348
g22093 and n22347_not n22348_not ; n22349
g22094 and n22346_not n22349 ; n22350
g22095 and n6219 n8365 ; n22351
g22096 and n22350 n22351_not ; n22352
g22097 and a[50] n22352_not ; n22353
g22098 and a[50] n22353_not ; n22354
g22099 and n22352_not n22353_not ; n22355
g22100 and n22354_not n22355_not ; n22356
g22101 and n22345_not n22356 ; n22357
g22102 and n22345 n22356_not ; n22358
g22103 and n22357_not n22358_not ; n22359
g22104 and n22265_not n22359_not ; n22360
g22105 and n22265 n22359 ; n22361
g22106 and n22360_not n22361_not ; n22362
g22107 and n22264_not n22362 ; n22363
g22108 and n22264 n22362_not ; n22364
g22109 and n22363_not n22364_not ; n22365
g22110 and n22253_not n22365 ; n22366
g22111 and n22253 n22365_not ; n22367
g22112 and n22366_not n22367_not ; n22368
g22113 and b[47] n6595 ; n22369
g22114 and b[45] n6902 ; n22370
g22115 and b[46] n6590 ; n22371
g22116 and n22370_not n22371_not ; n22372
g22117 and n22369_not n22372 ; n22373
g22118 and n6598 n7703 ; n22374
g22119 and n22373 n22374_not ; n22375
g22120 and a[44] n22375_not ; n22376
g22121 and a[44] n22376_not ; n22377
g22122 and n22375_not n22376_not ; n22378
g22123 and n22377_not n22378_not ; n22379
g22124 and n22368 n22379_not ; n22380
g22125 and n22368 n22380_not ; n22381
g22126 and n22379_not n22380_not ; n22382
g22127 and n22381_not n22382_not ; n22383
g22128 and n22078_not n22091_not ; n22384
g22129 and n22383 n22384 ; n22385
g22130 and n22383_not n22384_not ; n22386
g22131 and n22385_not n22386_not ; n22387
g22132 and b[50] n5777 ; n22388
g22133 and b[48] n6059 ; n22389
g22134 and b[49] n5772 ; n22390
g22135 and n22389_not n22390_not ; n22391
g22136 and n22388_not n22391 ; n22392
g22137 and n5780 n8949 ; n22393
g22138 and n22392 n22393_not ; n22394
g22139 and a[41] n22394_not ; n22395
g22140 and a[41] n22395_not ; n22396
g22141 and n22394_not n22395_not ; n22397
g22142 and n22396_not n22397_not ; n22398
g22143 and n22387_not n22398 ; n22399
g22144 and n22387 n22398_not ; n22400
g22145 and n22399_not n22400_not ; n22401
g22146 and n22252_not n22401 ; n22402
g22147 and n22252_not n22402_not ; n22403
g22148 and n22401 n22402_not ; n22404
g22149 and n22403_not n22404_not ; n22405
g22150 and n22251_not n22405_not ; n22406
g22151 and n22251 n22404_not ; n22407
g22152 and n22403_not n22407 ; n22408
g22153 and n22406_not n22408_not ; n22409
g22154 and n22240_not n22409 ; n22410
g22155 and n22240 n22409_not ; n22411
g22156 and n22410_not n22411_not ; n22412
g22157 and n22239_not n22412 ; n22413
g22158 and n22239_not n22413_not ; n22414
g22159 and n22412 n22413_not ; n22415
g22160 and n22414_not n22415_not ; n22416
g22161 and n22228 n22416_not ; n22417
g22162 and n22228 n22417_not ; n22418
g22163 and n22416_not n22417_not ; n22419
g22164 and n22418_not n22419_not ; n22420
g22165 and n22212_not n22420 ; n22421
g22166 and n22212 n22420_not ; n22422
g22167 and n22421_not n22422_not ; n22423
g22168 and n22197_not n22423 ; n22424
g22169 and n22197 n22423_not ; n22425
g22170 and n22424_not n22425_not ; n22426
g22171 and n22185_not n22426 ; n22427
g22172 and n22185 n22426_not ; n22428
g22173 and n22427_not n22428_not ; n22429
g22174 and n22184_not n22429 ; n22430
g22175 and n22184 n22429_not ; n22431
g22176 and n22430_not n22431_not ; f[89]
g22177 and n22194_not n22424_not ; n22433
g22178 and n22211_not n22422_not ; n22434
g22179 and b[63] n3050 ; n22435
g22180 and b[61] n3243 ; n22436
g22181 and b[62] n3045 ; n22437
g22182 and n22436_not n22437_not ; n22438
g22183 and n22435_not n22438 ; n22439
g22184 and n3053 n13771 ; n22440
g22185 and n22439 n22440_not ; n22441
g22186 and a[29] n22441_not ; n22442
g22187 and a[29] n22442_not ; n22443
g22188 and n22441_not n22442_not ; n22444
g22189 and n22443_not n22444_not ; n22445
g22190 and n22434_not n22445_not ; n22446
g22191 and n22434_not n22446_not ; n22447
g22192 and n22445_not n22446_not ; n22448
g22193 and n22447_not n22448_not ; n22449
g22194 and b[57] n4287 ; n22450
g22195 and b[55] n4532 ; n22451
g22196 and b[56] n4282 ; n22452
g22197 and n22451_not n22452_not ; n22453
g22198 and n22450_not n22453 ; n22454
g22199 and n4290 n11410 ; n22455
g22200 and n22454 n22455_not ; n22456
g22201 and a[35] n22456_not ; n22457
g22202 and a[35] n22457_not ; n22458
g22203 and n22456_not n22457_not ; n22459
g22204 and n22458_not n22459_not ; n22460
g22205 and n22402_not n22406_not ; n22461
g22206 and n22386_not n22400_not ; n22462
g22207 and n22360_not n22363_not ; n22463
g22208 and n22345_not n22356_not ; n22464
g22209 and n22342_not n22464_not ; n22465
g22210 and b[33] n11531 ; n22466
g22211 and b[31] n11896 ; n22467
g22212 and b[32] n11526 ; n22468
g22213 and n22467_not n22468_not ; n22469
g22214 and n22466_not n22469 ; n22470
g22215 and n4223 n11534 ; n22471
g22216 and n22470 n22471_not ; n22472
g22217 and a[59] n22472_not ; n22473
g22218 and a[59] n22473_not ; n22474
g22219 and n22472_not n22473_not ; n22475
g22220 and n22474_not n22475_not ; n22476
g22221 and n22311_not n22314_not ; n22477
g22222 and n22476 n22477 ; n22478
g22223 and n22476_not n22477_not ; n22479
g22224 and n22478_not n22479_not ; n22480
g22225 and n22294_not n22308_not ; n22481
g22226 and b[26] n13903 ; n22482
g22227 and b[27] n13488_not ; n22483
g22228 and n22482_not n22483_not ; n22484
g22229 and a[26]_not n22484_not ; n22485
g22230 and a[26] n22484 ; n22486
g22231 and n22485_not n22486_not ; n22487
g22232 and n22293_not n22487 ; n22488
g22233 and n22293 n22487_not ; n22489
g22234 and n22488_not n22489_not ; n22490
g22235 and n22481_not n22490 ; n22491
g22236 and n22481 n22490_not ; n22492
g22237 and n22491_not n22492_not ; n22493
g22238 and b[30] n12668 ; n22494
g22239 and b[28] n13047 ; n22495
g22240 and b[29] n12663 ; n22496
g22241 and n22495_not n22496_not ; n22497
g22242 and n22494_not n22497 ; n22498
g22243 and n3577 n12671 ; n22499
g22244 and n22498 n22499_not ; n22500
g22245 and a[62] n22500_not ; n22501
g22246 and a[62] n22501_not ; n22502
g22247 and n22500_not n22501_not ; n22503
g22248 and n22502_not n22503_not ; n22504
g22249 and n22493 n22504_not ; n22505
g22250 and n22493 n22505_not ; n22506
g22251 and n22504_not n22505_not ; n22507
g22252 and n22506_not n22507_not ; n22508
g22253 and n22480_not n22508 ; n22509
g22254 and n22480 n22508_not ; n22510
g22255 and n22509_not n22510_not ; n22511
g22256 and b[36] n10426 ; n22512
g22257 and b[34] n10796 ; n22513
g22258 and b[35] n10421 ; n22514
g22259 and n22513_not n22514_not ; n22515
g22260 and n22512_not n22515 ; n22516
g22261 and n4922 n10429 ; n22517
g22262 and n22516 n22517_not ; n22518
g22263 and a[56] n22518_not ; n22519
g22264 and a[56] n22519_not ; n22520
g22265 and n22518_not n22519_not ; n22521
g22266 and n22520_not n22521_not ; n22522
g22267 and n22511 n22522_not ; n22523
g22268 and n22511 n22523_not ; n22524
g22269 and n22522_not n22523_not ; n22525
g22270 and n22524_not n22525_not ; n22526
g22271 and n22317_not n22320_not ; n22527
g22272 and n22526 n22527 ; n22528
g22273 and n22526_not n22527_not ; n22529
g22274 and n22528_not n22529_not ; n22530
g22275 and b[39] n9339 ; n22531
g22276 and b[37] n9732 ; n22532
g22277 and b[38] n9334 ; n22533
g22278 and n22532_not n22533_not ; n22534
g22279 and n22531_not n22534 ; n22535
g22280 and n5451 n9342 ; n22536
g22281 and n22535 n22536_not ; n22537
g22282 and a[53] n22537_not ; n22538
g22283 and a[53] n22538_not ; n22539
g22284 and n22537_not n22538_not ; n22540
g22285 and n22539_not n22540_not ; n22541
g22286 and n22530 n22541_not ; n22542
g22287 and n22530 n22542_not ; n22543
g22288 and n22541_not n22542_not ; n22544
g22289 and n22543_not n22544_not ; n22545
g22290 and n22323_not n22337_not ; n22546
g22291 and n22545 n22546 ; n22547
g22292 and n22545_not n22546_not ; n22548
g22293 and n22547_not n22548_not ; n22549
g22294 and b[42] n8362 ; n22550
g22295 and b[40] n8715 ; n22551
g22296 and b[41] n8357 ; n22552
g22297 and n22551_not n22552_not ; n22553
g22298 and n22550_not n22553 ; n22554
g22299 and n6489 n8365 ; n22555
g22300 and n22554 n22555_not ; n22556
g22301 and a[50] n22556_not ; n22557
g22302 and a[50] n22557_not ; n22558
g22303 and n22556_not n22557_not ; n22559
g22304 and n22558_not n22559_not ; n22560
g22305 and n22549 n22560_not ; n22561
g22306 and n22549 n22561_not ; n22562
g22307 and n22560_not n22561_not ; n22563
g22308 and n22562_not n22563_not ; n22564
g22309 and n22465_not n22564 ; n22565
g22310 and n22465 n22564_not ; n22566
g22311 and n22565_not n22566_not ; n22567
g22312 and b[45] n7446 ; n22568
g22313 and b[43] n7787 ; n22569
g22314 and b[44] n7441 ; n22570
g22315 and n22569_not n22570_not ; n22571
g22316 and n22568_not n22571 ; n22572
g22317 and n7361 n7449 ; n22573
g22318 and n22572 n22573_not ; n22574
g22319 and a[47] n22574_not ; n22575
g22320 and a[47] n22575_not ; n22576
g22321 and n22574_not n22575_not ; n22577
g22322 and n22576_not n22577_not ; n22578
g22323 and n22567_not n22578_not ; n22579
g22324 and n22567 n22578 ; n22580
g22325 and n22579_not n22580_not ; n22581
g22326 and n22463 n22581_not ; n22582
g22327 and n22463_not n22581 ; n22583
g22328 and n22582_not n22583_not ; n22584
g22329 and b[48] n6595 ; n22585
g22330 and b[46] n6902 ; n22586
g22331 and b[47] n6590 ; n22587
g22332 and n22586_not n22587_not ; n22588
g22333 and n22585_not n22588 ; n22589
g22334 and n6598 n8009 ; n22590
g22335 and n22589 n22590_not ; n22591
g22336 and a[44] n22591_not ; n22592
g22337 and a[44] n22592_not ; n22593
g22338 and n22591_not n22592_not ; n22594
g22339 and n22593_not n22594_not ; n22595
g22340 and n22584 n22595_not ; n22596
g22341 and n22584 n22596_not ; n22597
g22342 and n22595_not n22596_not ; n22598
g22343 and n22597_not n22598_not ; n22599
g22344 and n22366_not n22380_not ; n22600
g22345 and n22599 n22600 ; n22601
g22346 and n22599_not n22600_not ; n22602
g22347 and n22601_not n22602_not ; n22603
g22348 and b[51] n5777 ; n22604
g22349 and b[49] n6059 ; n22605
g22350 and b[50] n5772 ; n22606
g22351 and n22605_not n22606_not ; n22607
g22352 and n22604_not n22607 ; n22608
g22353 and n5780 n8976 ; n22609
g22354 and n22608 n22609_not ; n22610
g22355 and a[41] n22610_not ; n22611
g22356 and a[41] n22611_not ; n22612
g22357 and n22610_not n22611_not ; n22613
g22358 and n22612_not n22613_not ; n22614
g22359 and n22603 n22614_not ; n22615
g22360 and n22603_not n22614 ; n22616
g22361 and n22462_not n22616_not ; n22617
g22362 and n22615_not n22617 ; n22618
g22363 and n22462_not n22618_not ; n22619
g22364 and n22615_not n22618_not ; n22620
g22365 and n22616_not n22620 ; n22621
g22366 and n22619_not n22621_not ; n22622
g22367 and b[54] n5035 ; n22623
g22368 and b[52] n5277 ; n22624
g22369 and b[53] n5030 ; n22625
g22370 and n22624_not n22625_not ; n22626
g22371 and n22623_not n22626 ; n22627
g22372 and n5038 n9998 ; n22628
g22373 and n22627 n22628_not ; n22629
g22374 and a[38] n22629_not ; n22630
g22375 and a[38] n22630_not ; n22631
g22376 and n22629_not n22630_not ; n22632
g22377 and n22631_not n22632_not ; n22633
g22378 and n22622 n22633 ; n22634
g22379 and n22622_not n22633_not ; n22635
g22380 and n22634_not n22635_not ; n22636
g22381 and n22461_not n22636 ; n22637
g22382 and n22461 n22636_not ; n22638
g22383 and n22637_not n22638_not ; n22639
g22384 and n22460_not n22639 ; n22640
g22385 and n22639 n22640_not ; n22641
g22386 and n22460_not n22640_not ; n22642
g22387 and n22641_not n22642_not ; n22643
g22388 and n22410_not n22413_not ; n22644
g22389 and n22643 n22644 ; n22645
g22390 and n22643_not n22644_not ; n22646
g22391 and n22645_not n22646_not ; n22647
g22392 and b[60] n3638 ; n22648
g22393 and b[58] n3843 ; n22649
g22394 and b[59] n3633 ; n22650
g22395 and n22649_not n22650_not ; n22651
g22396 and n22648_not n22651 ; n22652
g22397 and n3641 n12211 ; n22653
g22398 and n22652 n22653_not ; n22654
g22399 and a[32] n22654_not ; n22655
g22400 and a[32] n22655_not ; n22656
g22401 and n22654_not n22655_not ; n22657
g22402 and n22656_not n22657_not ; n22658
g22403 and n22227_not n22417_not ; n22659
g22404 and n22658 n22659 ; n22660
g22405 and n22658_not n22659_not ; n22661
g22406 and n22660_not n22661_not ; n22662
g22407 and n22647 n22662_not ; n22663
g22408 and n22647_not n22662 ; n22664
g22409 and n22663_not n22664_not ; n22665
g22410 and n22449_not n22665_not ; n22666
g22411 and n22449 n22665 ; n22667
g22412 and n22666_not n22667_not ; n22668
g22413 and n22433 n22668_not ; n22669
g22414 and n22433_not n22668 ; n22670
g22415 and n22669_not n22670_not ; n22671
g22416 and n22427_not n22430_not ; n22672
g22417 and n22671 n22672_not ; n22673
g22418 and n22671_not n22672 ; n22674
g22419 and n22673_not n22674_not ; f[90]
g22420 and n22647 n22662 ; n22676
g22421 and n22661_not n22676_not ; n22677
g22422 and b[62] n3243 ; n22678
g22423 and b[63] n3045 ; n22679
g22424 and n22678_not n22679_not ; n22680
g22425 and n3053_not n22680 ; n22681
g22426 and n13800 n22680 ; n22682
g22427 and n22681_not n22682_not ; n22683
g22428 and a[29] n22683_not ; n22684
g22429 and a[29]_not n22683 ; n22685
g22430 and n22684_not n22685_not ; n22686
g22431 and n22677_not n22686_not ; n22687
g22432 and n22677 n22686 ; n22688
g22433 and n22687_not n22688_not ; n22689
g22434 and b[61] n3638 ; n22690
g22435 and b[59] n3843 ; n22691
g22436 and b[60] n3633 ; n22692
g22437 and n22691_not n22692_not ; n22693
g22438 and n22690_not n22693 ; n22694
g22439 and n3641 n12969 ; n22695
g22440 and n22694 n22695_not ; n22696
g22441 and a[32] n22696_not ; n22697
g22442 and a[32] n22697_not ; n22698
g22443 and n22696_not n22697_not ; n22699
g22444 and n22698_not n22699_not ; n22700
g22445 and n22640_not n22646_not ; n22701
g22446 and n22700 n22701 ; n22702
g22447 and n22700_not n22701_not ; n22703
g22448 and n22702_not n22703_not ; n22704
g22449 and b[58] n4287 ; n22705
g22450 and b[56] n4532 ; n22706
g22451 and b[57] n4282 ; n22707
g22452 and n22706_not n22707_not ; n22708
g22453 and n22705_not n22708 ; n22709
g22454 and n4290 n11436 ; n22710
g22455 and n22709 n22710_not ; n22711
g22456 and a[35] n22711_not ; n22712
g22457 and a[35] n22712_not ; n22713
g22458 and n22711_not n22712_not ; n22714
g22459 and n22713_not n22714_not ; n22715
g22460 and n22635_not n22637_not ; n22716
g22461 and b[43] n8362 ; n22717
g22462 and b[41] n8715 ; n22718
g22463 and b[42] n8357 ; n22719
g22464 and n22718_not n22719_not ; n22720
g22465 and n22717_not n22720 ; n22721
g22466 and n6515 n8365 ; n22722
g22467 and n22721 n22722_not ; n22723
g22468 and a[50] n22723_not ; n22724
g22469 and a[50] n22724_not ; n22725
g22470 and n22723_not n22724_not ; n22726
g22471 and n22725_not n22726_not ; n22727
g22472 and n22542_not n22548_not ; n22728
g22473 and b[40] n9339 ; n22729
g22474 and b[38] n9732 ; n22730
g22475 and b[39] n9334 ; n22731
g22476 and n22730_not n22731_not ; n22732
g22477 and n22729_not n22732 ; n22733
g22478 and n5955 n9342 ; n22734
g22479 and n22733 n22734_not ; n22735
g22480 and a[53] n22735_not ; n22736
g22481 and a[53] n22736_not ; n22737
g22482 and n22735_not n22736_not ; n22738
g22483 and n22737_not n22738_not ; n22739
g22484 and n22523_not n22529_not ; n22740
g22485 and b[34] n11531 ; n22741
g22486 and b[32] n11896 ; n22742
g22487 and b[33] n11526 ; n22743
g22488 and n22742_not n22743_not ; n22744
g22489 and n22741_not n22744 ; n22745
g22490 and n4466 n11534 ; n22746
g22491 and n22745 n22746_not ; n22747
g22492 and a[59] n22747_not ; n22748
g22493 and a[59] n22748_not ; n22749
g22494 and n22747_not n22748_not ; n22750
g22495 and n22749_not n22750_not ; n22751
g22496 and b[27] n13903 ; n22752
g22497 and b[28] n13488_not ; n22753
g22498 and n22752_not n22753_not ; n22754
g22499 and n22485_not n22488_not ; n22755
g22500 and n22754_not n22755 ; n22756
g22501 and n22754 n22755_not ; n22757
g22502 and n22756_not n22757_not ; n22758
g22503 and b[31] n12668 ; n22759
g22504 and b[29] n13047 ; n22760
g22505 and b[30] n12663 ; n22761
g22506 and n22760_not n22761_not ; n22762
g22507 and n22759_not n22762 ; n22763
g22508 and n3796 n12671 ; n22764
g22509 and n22763 n22764_not ; n22765
g22510 and a[62] n22765_not ; n22766
g22511 and a[62] n22766_not ; n22767
g22512 and n22765_not n22766_not ; n22768
g22513 and n22767_not n22768_not ; n22769
g22514 and n22758_not n22769 ; n22770
g22515 and n22758 n22769_not ; n22771
g22516 and n22770_not n22771_not ; n22772
g22517 and n22491_not n22505_not ; n22773
g22518 and n22772 n22773_not ; n22774
g22519 and n22772_not n22773 ; n22775
g22520 and n22774_not n22775_not ; n22776
g22521 and n22751_not n22776 ; n22777
g22522 and n22776 n22777_not ; n22778
g22523 and n22751_not n22777_not ; n22779
g22524 and n22778_not n22779_not ; n22780
g22525 and n22479_not n22510_not ; n22781
g22526 and n22780_not n22781_not ; n22782
g22527 and n22780_not n22782_not ; n22783
g22528 and n22781_not n22782_not ; n22784
g22529 and n22783_not n22784_not ; n22785
g22530 and b[37] n10426 ; n22786
g22531 and b[35] n10796 ; n22787
g22532 and b[36] n10421 ; n22788
g22533 and n22787_not n22788_not ; n22789
g22534 and n22786_not n22789 ; n22790
g22535 and n5181 n10429 ; n22791
g22536 and n22790 n22791_not ; n22792
g22537 and a[56] n22792_not ; n22793
g22538 and a[56] n22793_not ; n22794
g22539 and n22792_not n22793_not ; n22795
g22540 and n22794_not n22795_not ; n22796
g22541 and n22785_not n22796 ; n22797
g22542 and n22785 n22796_not ; n22798
g22543 and n22797_not n22798_not ; n22799
g22544 and n22740_not n22799_not ; n22800
g22545 and n22740_not n22800_not ; n22801
g22546 and n22799_not n22800_not ; n22802
g22547 and n22801_not n22802_not ; n22803
g22548 and n22739_not n22803_not ; n22804
g22549 and n22739 n22802_not ; n22805
g22550 and n22801_not n22805 ; n22806
g22551 and n22804_not n22806_not ; n22807
g22552 and n22728_not n22807 ; n22808
g22553 and n22728 n22807_not ; n22809
g22554 and n22808_not n22809_not ; n22810
g22555 and n22727_not n22810 ; n22811
g22556 and n22810 n22811_not ; n22812
g22557 and n22727_not n22811_not ; n22813
g22558 and n22812_not n22813_not ; n22814
g22559 and n22465_not n22564_not ; n22815
g22560 and n22561_not n22815_not ; n22816
g22561 and n22814 n22816 ; n22817
g22562 and n22814_not n22816_not ; n22818
g22563 and n22817_not n22818_not ; n22819
g22564 and b[46] n7446 ; n22820
g22565 and b[44] n7787 ; n22821
g22566 and b[45] n7441 ; n22822
g22567 and n22821_not n22822_not ; n22823
g22568 and n22820_not n22823 ; n22824
g22569 and n7449 n7677 ; n22825
g22570 and n22824 n22825_not ; n22826
g22571 and a[47] n22826_not ; n22827
g22572 and a[47] n22827_not ; n22828
g22573 and n22826_not n22827_not ; n22829
g22574 and n22828_not n22829_not ; n22830
g22575 and n22819 n22830_not ; n22831
g22576 and n22819 n22831_not ; n22832
g22577 and n22830_not n22831_not ; n22833
g22578 and n22832_not n22833_not ; n22834
g22579 and n22579_not n22583_not ; n22835
g22580 and n22834 n22835 ; n22836
g22581 and n22834_not n22835_not ; n22837
g22582 and n22836_not n22837_not ; n22838
g22583 and b[49] n6595 ; n22839
g22584 and b[47] n6902 ; n22840
g22585 and b[48] n6590 ; n22841
g22586 and n22840_not n22841_not ; n22842
g22587 and n22839_not n22842 ; n22843
g22588 and n6598 n8625 ; n22844
g22589 and n22843 n22844_not ; n22845
g22590 and a[44] n22845_not ; n22846
g22591 and a[44] n22846_not ; n22847
g22592 and n22845_not n22846_not ; n22848
g22593 and n22847_not n22848_not ; n22849
g22594 and n22838 n22849_not ; n22850
g22595 and n22838 n22850_not ; n22851
g22596 and n22849_not n22850_not ; n22852
g22597 and n22851_not n22852_not ; n22853
g22598 and n22596_not n22602_not ; n22854
g22599 and n22853 n22854 ; n22855
g22600 and n22853_not n22854_not ; n22856
g22601 and n22855_not n22856_not ; n22857
g22602 and b[52] n5777 ; n22858
g22603 and b[50] n6059 ; n22859
g22604 and b[51] n5772 ; n22860
g22605 and n22859_not n22860_not ; n22861
g22606 and n22858_not n22861 ; n22862
g22607 and n5780 n9628 ; n22863
g22608 and n22862 n22863_not ; n22864
g22609 and a[41] n22864_not ; n22865
g22610 and a[41] n22865_not ; n22866
g22611 and n22864_not n22865_not ; n22867
g22612 and n22866_not n22867_not ; n22868
g22613 and n22857 n22868_not ; n22869
g22614 and n22857 n22869_not ; n22870
g22615 and n22868_not n22869_not ; n22871
g22616 and n22870_not n22871_not ; n22872
g22617 and n22620_not n22872 ; n22873
g22618 and n22620 n22872_not ; n22874
g22619 and n22873_not n22874_not ; n22875
g22620 and b[55] n5035 ; n22876
g22621 and b[53] n5277 ; n22877
g22622 and b[54] n5030 ; n22878
g22623 and n22877_not n22878_not ; n22879
g22624 and n22876_not n22879 ; n22880
g22625 and n5038 n10684 ; n22881
g22626 and n22880 n22881_not ; n22882
g22627 and a[38] n22882_not ; n22883
g22628 and a[38] n22883_not ; n22884
g22629 and n22882_not n22883_not ; n22885
g22630 and n22884_not n22885_not ; n22886
g22631 and n22875_not n22886_not ; n22887
g22632 and n22875 n22886 ; n22888
g22633 and n22887_not n22888_not ; n22889
g22634 and n22716_not n22889 ; n22890
g22635 and n22716 n22889_not ; n22891
g22636 and n22890_not n22891_not ; n22892
g22637 and n22715_not n22892 ; n22893
g22638 and n22892 n22893_not ; n22894
g22639 and n22715_not n22893_not ; n22895
g22640 and n22894_not n22895_not ; n22896
g22641 and n22704 n22896_not ; n22897
g22642 and n22704_not n22896 ; n22898
g22643 and n22689 n22898_not ; n22899
g22644 and n22897_not n22899 ; n22900
g22645 and n22689 n22900_not ; n22901
g22646 and n22898_not n22900_not ; n22902
g22647 and n22897_not n22902 ; n22903
g22648 and n22901_not n22903_not ; n22904
g22649 and n22446_not n22666_not ; n22905
g22650 and n22904 n22905 ; n22906
g22651 and n22904_not n22905_not ; n22907
g22652 and n22906_not n22907_not ; n22908
g22653 and n22670_not n22673_not ; n22909
g22654 and n22908 n22909_not ; n22910
g22655 and n22908_not n22909 ; n22911
g22656 and n22910_not n22911_not ; f[91]
g22657 and n22907_not n22910_not ; n22913
g22658 and n22687_not n22900_not ; n22914
g22659 and n22703_not n22897_not ; n22915
g22660 and b[63] n3243 ; n22916
g22661 and n3053 n13797 ; n22917
g22662 and n22916_not n22917_not ; n22918
g22663 and a[29] n22918_not ; n22919
g22664 and a[29] n22919_not ; n22920
g22665 and n22918_not n22919_not ; n22921
g22666 and n22920_not n22921_not ; n22922
g22667 and n22915_not n22922_not ; n22923
g22668 and n22915_not n22923_not ; n22924
g22669 and n22922_not n22923_not ; n22925
g22670 and n22924_not n22925_not ; n22926
g22671 and b[62] n3638 ; n22927
g22672 and b[60] n3843 ; n22928
g22673 and b[61] n3633 ; n22929
g22674 and n22928_not n22929_not ; n22930
g22675 and n22927_not n22930 ; n22931
g22676 and n3641 n13370 ; n22932
g22677 and n22931 n22932_not ; n22933
g22678 and a[32] n22933_not ; n22934
g22679 and a[32] n22934_not ; n22935
g22680 and n22933_not n22934_not ; n22936
g22681 and n22935_not n22936_not ; n22937
g22682 and n22890_not n22893_not ; n22938
g22683 and n22937 n22938 ; n22939
g22684 and n22937_not n22938_not ; n22940
g22685 and n22939_not n22940_not ; n22941
g22686 and n22620_not n22872_not ; n22942
g22687 and n22887_not n22942_not ; n22943
g22688 and b[56] n5035 ; n22944
g22689 and b[54] n5277 ; n22945
g22690 and b[55] n5030 ; n22946
g22691 and n22945_not n22946_not ; n22947
g22692 and n22944_not n22947 ; n22948
g22693 and n5038 n10708 ; n22949
g22694 and n22948 n22949_not ; n22950
g22695 and a[38] n22950_not ; n22951
g22696 and a[38] n22951_not ; n22952
g22697 and n22950_not n22951_not ; n22953
g22698 and n22952_not n22953_not ; n22954
g22699 and n22856_not n22869_not ; n22955
g22700 and b[53] n5777 ; n22956
g22701 and b[51] n6059 ; n22957
g22702 and b[52] n5772 ; n22958
g22703 and n22957_not n22958_not ; n22959
g22704 and n22956_not n22959 ; n22960
g22705 and n5780 n9972 ; n22961
g22706 and n22960 n22961_not ; n22962
g22707 and a[41] n22962_not ; n22963
g22708 and a[41] n22963_not ; n22964
g22709 and n22962_not n22963_not ; n22965
g22710 and n22964_not n22965_not ; n22966
g22711 and n22837_not n22850_not ; n22967
g22712 and n22808_not n22811_not ; n22968
g22713 and b[44] n8362 ; n22969
g22714 and b[42] n8715 ; n22970
g22715 and b[43] n8357 ; n22971
g22716 and n22970_not n22971_not ; n22972
g22717 and n22969_not n22972 ; n22973
g22718 and n7072 n8365 ; n22974
g22719 and n22973 n22974_not ; n22975
g22720 and a[50] n22975_not ; n22976
g22721 and a[50] n22976_not ; n22977
g22722 and n22975_not n22976_not ; n22978
g22723 and n22977_not n22978_not ; n22979
g22724 and n22800_not n22804_not ; n22980
g22725 and n22774_not n22777_not ; n22981
g22726 and b[35] n11531 ; n22982
g22727 and b[33] n11896 ; n22983
g22728 and b[34] n11526 ; n22984
g22729 and n22983_not n22984_not ; n22985
g22730 and n22982_not n22985 ; n22986
g22731 and n4696 n11534 ; n22987
g22732 and n22986 n22987_not ; n22988
g22733 and a[59] n22988_not ; n22989
g22734 and a[59] n22989_not ; n22990
g22735 and n22988_not n22989_not ; n22991
g22736 and n22990_not n22991_not ; n22992
g22737 and n22757_not n22771_not ; n22993
g22738 and b[28] n13903 ; n22994
g22739 and b[29] n13488_not ; n22995
g22740 and n22994_not n22995_not ; n22996
g22741 and n22754 n22996_not ; n22997
g22742 and n22754_not n22996 ; n22998
g22743 and n22993_not n22998_not ; n22999
g22744 and n22997_not n22999 ; n23000
g22745 and n22993_not n23000_not ; n23001
g22746 and n22998_not n23000_not ; n23002
g22747 and n22997_not n23002 ; n23003
g22748 and n23001_not n23003_not ; n23004
g22749 and b[32] n12668 ; n23005
g22750 and b[30] n13047 ; n23006
g22751 and b[31] n12663 ; n23007
g22752 and n23006_not n23007_not ; n23008
g22753 and n23005_not n23008 ; n23009
g22754 and n4013 n12671 ; n23010
g22755 and n23009 n23010_not ; n23011
g22756 and a[62] n23011_not ; n23012
g22757 and a[62] n23012_not ; n23013
g22758 and n23011_not n23012_not ; n23014
g22759 and n23013_not n23014_not ; n23015
g22760 and n23004_not n23015 ; n23016
g22761 and n23004 n23015_not ; n23017
g22762 and n23016_not n23017_not ; n23018
g22763 and n22992_not n23018_not ; n23019
g22764 and n22992 n23018 ; n23020
g22765 and n23019_not n23020_not ; n23021
g22766 and n22981_not n23021 ; n23022
g22767 and n22981 n23021_not ; n23023
g22768 and n23022_not n23023_not ; n23024
g22769 and b[38] n10426 ; n23025
g22770 and b[36] n10796 ; n23026
g22771 and b[37] n10421 ; n23027
g22772 and n23026_not n23027_not ; n23028
g22773 and n23025_not n23028 ; n23029
g22774 and n5205 n10429 ; n23030
g22775 and n23029 n23030_not ; n23031
g22776 and a[56] n23031_not ; n23032
g22777 and a[56] n23032_not ; n23033
g22778 and n23031_not n23032_not ; n23034
g22779 and n23033_not n23034_not ; n23035
g22780 and n23024 n23035_not ; n23036
g22781 and n23024 n23036_not ; n23037
g22782 and n23035_not n23036_not ; n23038
g22783 and n23037_not n23038_not ; n23039
g22784 and n22785_not n22796_not ; n23040
g22785 and n22782_not n23040_not ; n23041
g22786 and n23039_not n23041_not ; n23042
g22787 and n23039_not n23042_not ; n23043
g22788 and n23041_not n23042_not ; n23044
g22789 and n23043_not n23044_not ; n23045
g22790 and b[41] n9339 ; n23046
g22791 and b[39] n9732 ; n23047
g22792 and b[40] n9334 ; n23048
g22793 and n23047_not n23048_not ; n23049
g22794 and n23046_not n23049 ; n23050
g22795 and n6219 n9342 ; n23051
g22796 and n23050 n23051_not ; n23052
g22797 and a[53] n23052_not ; n23053
g22798 and a[53] n23053_not ; n23054
g22799 and n23052_not n23053_not ; n23055
g22800 and n23054_not n23055_not ; n23056
g22801 and n23045_not n23056 ; n23057
g22802 and n23045 n23056_not ; n23058
g22803 and n23057_not n23058_not ; n23059
g22804 and n22980_not n23059_not ; n23060
g22805 and n22980 n23059 ; n23061
g22806 and n23060_not n23061_not ; n23062
g22807 and n22979_not n23062 ; n23063
g22808 and n22979 n23062_not ; n23064
g22809 and n23063_not n23064_not ; n23065
g22810 and n22968_not n23065 ; n23066
g22811 and n22968 n23065_not ; n23067
g22812 and n23066_not n23067_not ; n23068
g22813 and b[47] n7446 ; n23069
g22814 and b[45] n7787 ; n23070
g22815 and b[46] n7441 ; n23071
g22816 and n23070_not n23071_not ; n23072
g22817 and n23069_not n23072 ; n23073
g22818 and n7449 n7703 ; n23074
g22819 and n23073 n23074_not ; n23075
g22820 and a[47] n23075_not ; n23076
g22821 and a[47] n23076_not ; n23077
g22822 and n23075_not n23076_not ; n23078
g22823 and n23077_not n23078_not ; n23079
g22824 and n23068 n23079_not ; n23080
g22825 and n23068 n23080_not ; n23081
g22826 and n23079_not n23080_not ; n23082
g22827 and n23081_not n23082_not ; n23083
g22828 and n22818_not n22831_not ; n23084
g22829 and n23083 n23084 ; n23085
g22830 and n23083_not n23084_not ; n23086
g22831 and n23085_not n23086_not ; n23087
g22832 and b[50] n6595 ; n23088
g22833 and b[48] n6902 ; n23089
g22834 and b[49] n6590 ; n23090
g22835 and n23089_not n23090_not ; n23091
g22836 and n23088_not n23091 ; n23092
g22837 and n6598 n8949 ; n23093
g22838 and n23092 n23093_not ; n23094
g22839 and a[44] n23094_not ; n23095
g22840 and a[44] n23095_not ; n23096
g22841 and n23094_not n23095_not ; n23097
g22842 and n23096_not n23097_not ; n23098
g22843 and n23087_not n23098 ; n23099
g22844 and n23087 n23098_not ; n23100
g22845 and n23099_not n23100_not ; n23101
g22846 and n22967_not n23101 ; n23102
g22847 and n22967_not n23102_not ; n23103
g22848 and n23101 n23102_not ; n23104
g22849 and n23103_not n23104_not ; n23105
g22850 and n22966_not n23105_not ; n23106
g22851 and n22966 n23104_not ; n23107
g22852 and n23103_not n23107 ; n23108
g22853 and n23106_not n23108_not ; n23109
g22854 and n22955_not n23109 ; n23110
g22855 and n22955 n23109_not ; n23111
g22856 and n23110_not n23111_not ; n23112
g22857 and n22954_not n23112 ; n23113
g22858 and n22954 n23112_not ; n23114
g22859 and n23113_not n23114_not ; n23115
g22860 and n22943_not n23115 ; n23116
g22861 and n22943 n23115_not ; n23117
g22862 and n23116_not n23117_not ; n23118
g22863 and b[59] n4287 ; n23119
g22864 and b[57] n4532 ; n23120
g22865 and b[58] n4282 ; n23121
g22866 and n23120_not n23121_not ; n23122
g22867 and n23119_not n23122 ; n23123
g22868 and n4290 n12179 ; n23124
g22869 and n23123 n23124_not ; n23125
g22870 and a[35] n23125_not ; n23126
g22871 and a[35] n23126_not ; n23127
g22872 and n23125_not n23126_not ; n23128
g22873 and n23127_not n23128_not ; n23129
g22874 and n23118 n23129_not ; n23130
g22875 and n23118 n23130_not ; n23131
g22876 and n23129_not n23130_not ; n23132
g22877 and n23131_not n23132_not ; n23133
g22878 and n22941_not n23133 ; n23134
g22879 and n22941 n23133_not ; n23135
g22880 and n23134_not n23135_not ; n23136
g22881 and n22926_not n23136 ; n23137
g22882 and n22926 n23136_not ; n23138
g22883 and n23137_not n23138_not ; n23139
g22884 and n22914_not n23139 ; n23140
g22885 and n22914_not n23140_not ; n23141
g22886 and n23139 n23140_not ; n23142
g22887 and n23141_not n23142_not ; n23143
g22888 and n22913_not n23143_not ; n23144
g22889 and n22913 n23142_not ; n23145
g22890 and n23141_not n23145 ; n23146
g22891 and n23144_not n23146_not ; f[92]
g22892 and n23140_not n23144_not ; n23148
g22893 and n22923_not n23137_not ; n23149
g22894 and b[57] n5035 ; n23150
g22895 and b[55] n5277 ; n23151
g22896 and b[56] n5030 ; n23152
g22897 and n23151_not n23152_not ; n23153
g22898 and n23150_not n23153 ; n23154
g22899 and n5038 n11410 ; n23155
g22900 and n23154 n23155_not ; n23156
g22901 and a[38] n23156_not ; n23157
g22902 and a[38] n23157_not ; n23158
g22903 and n23156_not n23157_not ; n23159
g22904 and n23158_not n23159_not ; n23160
g22905 and n23102_not n23106_not ; n23161
g22906 and n23086_not n23100_not ; n23162
g22907 and n23060_not n23063_not ; n23163
g22908 and n23045_not n23056_not ; n23164
g22909 and n23042_not n23164_not ; n23165
g22910 and b[39] n10426 ; n23166
g22911 and b[37] n10796 ; n23167
g22912 and b[38] n10421 ; n23168
g22913 and n23167_not n23168_not ; n23169
g22914 and n23166_not n23169 ; n23170
g22915 and n5451 n10429 ; n23171
g22916 and n23170 n23171_not ; n23172
g22917 and a[56] n23172_not ; n23173
g22918 and a[56] n23173_not ; n23174
g22919 and n23172_not n23173_not ; n23175
g22920 and n23174_not n23175_not ; n23176
g22921 and n23004_not n23015_not ; n23177
g22922 and n23019_not n23177_not ; n23178
g22923 and b[29] n13903 ; n23179
g22924 and b[30] n13488_not ; n23180
g22925 and n23179_not n23180_not ; n23181
g22926 and a[29]_not n23181_not ; n23182
g22927 and a[29] n23181 ; n23183
g22928 and n23182_not n23183_not ; n23184
g22929 and n22996_not n23184 ; n23185
g22930 and n22996_not n23185_not ; n23186
g22931 and n23184 n23185_not ; n23187
g22932 and n23186_not n23187_not ; n23188
g22933 and n23002_not n23188_not ; n23189
g22934 and n23002_not n23189_not ; n23190
g22935 and n23188_not n23189_not ; n23191
g22936 and n23190_not n23191_not ; n23192
g22937 and b[33] n12668 ; n23193
g22938 and b[31] n13047 ; n23194
g22939 and b[32] n12663 ; n23195
g22940 and n23194_not n23195_not ; n23196
g22941 and n23193_not n23196 ; n23197
g22942 and n4223 n12671 ; n23198
g22943 and n23197 n23198_not ; n23199
g22944 and a[62] n23199_not ; n23200
g22945 and a[62] n23200_not ; n23201
g22946 and n23199_not n23200_not ; n23202
g22947 and n23201_not n23202_not ; n23203
g22948 and n23192_not n23203 ; n23204
g22949 and n23192 n23203_not ; n23205
g22950 and n23204_not n23205_not ; n23206
g22951 and b[36] n11531 ; n23207
g22952 and b[34] n11896 ; n23208
g22953 and b[35] n11526 ; n23209
g22954 and n23208_not n23209_not ; n23210
g22955 and n23207_not n23210 ; n23211
g22956 and n4922 n11534 ; n23212
g22957 and n23211 n23212_not ; n23213
g22958 and a[59] n23213_not ; n23214
g22959 and a[59] n23214_not ; n23215
g22960 and n23213_not n23214_not ; n23216
g22961 and n23215_not n23216_not ; n23217
g22962 and n23206_not n23217_not ; n23218
g22963 and n23206 n23217 ; n23219
g22964 and n23218_not n23219_not ; n23220
g22965 and n23178_not n23220 ; n23221
g22966 and n23178 n23220_not ; n23222
g22967 and n23221_not n23222_not ; n23223
g22968 and n23176_not n23223 ; n23224
g22969 and n23223 n23224_not ; n23225
g22970 and n23176_not n23224_not ; n23226
g22971 and n23225_not n23226_not ; n23227
g22972 and n23022_not n23036_not ; n23228
g22973 and n23227 n23228 ; n23229
g22974 and n23227_not n23228_not ; n23230
g22975 and n23229_not n23230_not ; n23231
g22976 and b[42] n9339 ; n23232
g22977 and b[40] n9732 ; n23233
g22978 and b[41] n9334 ; n23234
g22979 and n23233_not n23234_not ; n23235
g22980 and n23232_not n23235 ; n23236
g22981 and n6489 n9342 ; n23237
g22982 and n23236 n23237_not ; n23238
g22983 and a[53] n23238_not ; n23239
g22984 and a[53] n23239_not ; n23240
g22985 and n23238_not n23239_not ; n23241
g22986 and n23240_not n23241_not ; n23242
g22987 and n23231 n23242_not ; n23243
g22988 and n23231 n23243_not ; n23244
g22989 and n23242_not n23243_not ; n23245
g22990 and n23244_not n23245_not ; n23246
g22991 and n23165_not n23246 ; n23247
g22992 and n23165 n23246_not ; n23248
g22993 and n23247_not n23248_not ; n23249
g22994 and b[45] n8362 ; n23250
g22995 and b[43] n8715 ; n23251
g22996 and b[44] n8357 ; n23252
g22997 and n23251_not n23252_not ; n23253
g22998 and n23250_not n23253 ; n23254
g22999 and n7361 n8365 ; n23255
g23000 and n23254 n23255_not ; n23256
g23001 and a[50] n23256_not ; n23257
g23002 and a[50] n23257_not ; n23258
g23003 and n23256_not n23257_not ; n23259
g23004 and n23258_not n23259_not ; n23260
g23005 and n23249_not n23260_not ; n23261
g23006 and n23249 n23260 ; n23262
g23007 and n23261_not n23262_not ; n23263
g23008 and n23163 n23263_not ; n23264
g23009 and n23163_not n23263 ; n23265
g23010 and n23264_not n23265_not ; n23266
g23011 and b[48] n7446 ; n23267
g23012 and b[46] n7787 ; n23268
g23013 and b[47] n7441 ; n23269
g23014 and n23268_not n23269_not ; n23270
g23015 and n23267_not n23270 ; n23271
g23016 and n7449 n8009 ; n23272
g23017 and n23271 n23272_not ; n23273
g23018 and a[47] n23273_not ; n23274
g23019 and a[47] n23274_not ; n23275
g23020 and n23273_not n23274_not ; n23276
g23021 and n23275_not n23276_not ; n23277
g23022 and n23266 n23277_not ; n23278
g23023 and n23266 n23278_not ; n23279
g23024 and n23277_not n23278_not ; n23280
g23025 and n23279_not n23280_not ; n23281
g23026 and n23066_not n23080_not ; n23282
g23027 and n23281 n23282 ; n23283
g23028 and n23281_not n23282_not ; n23284
g23029 and n23283_not n23284_not ; n23285
g23030 and b[51] n6595 ; n23286
g23031 and b[49] n6902 ; n23287
g23032 and b[50] n6590 ; n23288
g23033 and n23287_not n23288_not ; n23289
g23034 and n23286_not n23289 ; n23290
g23035 and n6598 n8976 ; n23291
g23036 and n23290 n23291_not ; n23292
g23037 and a[44] n23292_not ; n23293
g23038 and a[44] n23293_not ; n23294
g23039 and n23292_not n23293_not ; n23295
g23040 and n23294_not n23295_not ; n23296
g23041 and n23285 n23296_not ; n23297
g23042 and n23285_not n23296 ; n23298
g23043 and n23162_not n23298_not ; n23299
g23044 and n23297_not n23299 ; n23300
g23045 and n23162_not n23300_not ; n23301
g23046 and n23297_not n23300_not ; n23302
g23047 and n23298_not n23302 ; n23303
g23048 and n23301_not n23303_not ; n23304
g23049 and b[54] n5777 ; n23305
g23050 and b[52] n6059 ; n23306
g23051 and b[53] n5772 ; n23307
g23052 and n23306_not n23307_not ; n23308
g23053 and n23305_not n23308 ; n23309
g23054 and n5780 n9998 ; n23310
g23055 and n23309 n23310_not ; n23311
g23056 and a[41] n23311_not ; n23312
g23057 and a[41] n23312_not ; n23313
g23058 and n23311_not n23312_not ; n23314
g23059 and n23313_not n23314_not ; n23315
g23060 and n23304 n23315 ; n23316
g23061 and n23304_not n23315_not ; n23317
g23062 and n23316_not n23317_not ; n23318
g23063 and n23161_not n23318 ; n23319
g23064 and n23161 n23318_not ; n23320
g23065 and n23319_not n23320_not ; n23321
g23066 and n23160_not n23321 ; n23322
g23067 and n23321 n23322_not ; n23323
g23068 and n23160_not n23322_not ; n23324
g23069 and n23323_not n23324_not ; n23325
g23070 and n23110_not n23113_not ; n23326
g23071 and n23325 n23326 ; n23327
g23072 and n23325_not n23326_not ; n23328
g23073 and n23327_not n23328_not ; n23329
g23074 and b[60] n4287 ; n23330
g23075 and b[58] n4532 ; n23331
g23076 and b[59] n4282 ; n23332
g23077 and n23331_not n23332_not ; n23333
g23078 and n23330_not n23333 ; n23334
g23079 and n4290 n12211 ; n23335
g23080 and n23334 n23335_not ; n23336
g23081 and a[35] n23336_not ; n23337
g23082 and a[35] n23337_not ; n23338
g23083 and n23336_not n23337_not ; n23339
g23084 and n23338_not n23339_not ; n23340
g23085 and n23329 n23340_not ; n23341
g23086 and n23329 n23341_not ; n23342
g23087 and n23340_not n23341_not ; n23343
g23088 and n23342_not n23343_not ; n23344
g23089 and n23116_not n23130_not ; n23345
g23090 and n23344 n23345 ; n23346
g23091 and n23344_not n23345_not ; n23347
g23092 and n23346_not n23347_not ; n23348
g23093 and n22940_not n23135_not ; n23349
g23094 and b[63] n3638 ; n23350
g23095 and b[61] n3843 ; n23351
g23096 and b[62] n3633 ; n23352
g23097 and n23351_not n23352_not ; n23353
g23098 and n23350_not n23353 ; n23354
g23099 and n3641 n13771 ; n23355
g23100 and n23354 n23355_not ; n23356
g23101 and a[32] n23356_not ; n23357
g23102 and a[32] n23357_not ; n23358
g23103 and n23356_not n23357_not ; n23359
g23104 and n23358_not n23359_not ; n23360
g23105 and n23349_not n23360_not ; n23361
g23106 and n23349_not n23361_not ; n23362
g23107 and n23360_not n23361_not ; n23363
g23108 and n23362_not n23363_not ; n23364
g23109 and n23348_not n23364 ; n23365
g23110 and n23348 n23364_not ; n23366
g23111 and n23365_not n23366_not ; n23367
g23112 and n23149_not n23367 ; n23368
g23113 and n23149 n23367_not ; n23369
g23114 and n23368_not n23369_not ; n23370
g23115 and n23148_not n23370 ; n23371
g23116 and n23148 n23370_not ; n23372
g23117 and n23371_not n23372_not ; f[93]
g23118 and n23341_not n23347_not ; n23374
g23119 and b[62] n3843 ; n23375
g23120 and b[63] n3633 ; n23376
g23121 and n23375_not n23376_not ; n23377
g23122 and n3641_not n23377 ; n23378
g23123 and n13800 n23377 ; n23379
g23124 and n23378_not n23379_not ; n23380
g23125 and a[32] n23380_not ; n23381
g23126 and a[32]_not n23380 ; n23382
g23127 and n23381_not n23382_not ; n23383
g23128 and n23374_not n23383_not ; n23384
g23129 and n23374 n23383 ; n23385
g23130 and n23384_not n23385_not ; n23386
g23131 and b[58] n5035 ; n23387
g23132 and b[56] n5277 ; n23388
g23133 and b[57] n5030 ; n23389
g23134 and n23388_not n23389_not ; n23390
g23135 and n23387_not n23390 ; n23391
g23136 and n5038 n11436 ; n23392
g23137 and n23391 n23392_not ; n23393
g23138 and a[38] n23393_not ; n23394
g23139 and a[38] n23394_not ; n23395
g23140 and n23393_not n23394_not ; n23396
g23141 and n23395_not n23396_not ; n23397
g23142 and n23317_not n23319_not ; n23398
g23143 and b[43] n9339 ; n23399
g23144 and b[41] n9732 ; n23400
g23145 and b[42] n9334 ; n23401
g23146 and n23400_not n23401_not ; n23402
g23147 and n23399_not n23402 ; n23403
g23148 and n6515 n9342 ; n23404
g23149 and n23403 n23404_not ; n23405
g23150 and a[53] n23405_not ; n23406
g23151 and a[53] n23406_not ; n23407
g23152 and n23405_not n23406_not ; n23408
g23153 and n23407_not n23408_not ; n23409
g23154 and n23224_not n23230_not ; n23410
g23155 and b[40] n10426 ; n23411
g23156 and b[38] n10796 ; n23412
g23157 and b[39] n10421 ; n23413
g23158 and n23412_not n23413_not ; n23414
g23159 and n23411_not n23414 ; n23415
g23160 and n5955 n10429 ; n23416
g23161 and n23415 n23416_not ; n23417
g23162 and a[56] n23417_not ; n23418
g23163 and a[56] n23418_not ; n23419
g23164 and n23417_not n23418_not ; n23420
g23165 and n23419_not n23420_not ; n23421
g23166 and n23218_not n23221_not ; n23422
g23167 and b[37] n11531 ; n23423
g23168 and b[35] n11896 ; n23424
g23169 and b[36] n11526 ; n23425
g23170 and n23424_not n23425_not ; n23426
g23171 and n23423_not n23426 ; n23427
g23172 and n5181 n11534 ; n23428
g23173 and n23427 n23428_not ; n23429
g23174 and a[59] n23429_not ; n23430
g23175 and a[59] n23430_not ; n23431
g23176 and n23429_not n23430_not ; n23432
g23177 and n23431_not n23432_not ; n23433
g23178 and n23192_not n23203_not ; n23434
g23179 and n23189_not n23434_not ; n23435
g23180 and b[30] n13903 ; n23436
g23181 and b[31] n13488_not ; n23437
g23182 and n23436_not n23437_not ; n23438
g23183 and n23182_not n23185_not ; n23439
g23184 and n23438_not n23439 ; n23440
g23185 and n23438 n23439_not ; n23441
g23186 and n23440_not n23441_not ; n23442
g23187 and b[34] n12668 ; n23443
g23188 and b[32] n13047 ; n23444
g23189 and b[33] n12663 ; n23445
g23190 and n23444_not n23445_not ; n23446
g23191 and n23443_not n23446 ; n23447
g23192 and n4466 n12671 ; n23448
g23193 and n23447 n23448_not ; n23449
g23194 and a[62] n23449_not ; n23450
g23195 and a[62] n23450_not ; n23451
g23196 and n23449_not n23450_not ; n23452
g23197 and n23451_not n23452_not ; n23453
g23198 and n23442_not n23453 ; n23454
g23199 and n23442 n23453_not ; n23455
g23200 and n23454_not n23455_not ; n23456
g23201 and n23435_not n23456 ; n23457
g23202 and n23435_not n23457_not ; n23458
g23203 and n23456 n23457_not ; n23459
g23204 and n23458_not n23459_not ; n23460
g23205 and n23433_not n23460_not ; n23461
g23206 and n23433 n23459_not ; n23462
g23207 and n23458_not n23462 ; n23463
g23208 and n23461_not n23463_not ; n23464
g23209 and n23422_not n23464 ; n23465
g23210 and n23422_not n23465_not ; n23466
g23211 and n23464 n23465_not ; n23467
g23212 and n23466_not n23467_not ; n23468
g23213 and n23421_not n23468_not ; n23469
g23214 and n23421 n23467_not ; n23470
g23215 and n23466_not n23470 ; n23471
g23216 and n23469_not n23471_not ; n23472
g23217 and n23410_not n23472 ; n23473
g23218 and n23410 n23472_not ; n23474
g23219 and n23473_not n23474_not ; n23475
g23220 and n23409_not n23475 ; n23476
g23221 and n23475 n23476_not ; n23477
g23222 and n23409_not n23476_not ; n23478
g23223 and n23477_not n23478_not ; n23479
g23224 and n23165_not n23246_not ; n23480
g23225 and n23243_not n23480_not ; n23481
g23226 and n23479 n23481 ; n23482
g23227 and n23479_not n23481_not ; n23483
g23228 and n23482_not n23483_not ; n23484
g23229 and b[46] n8362 ; n23485
g23230 and b[44] n8715 ; n23486
g23231 and b[45] n8357 ; n23487
g23232 and n23486_not n23487_not ; n23488
g23233 and n23485_not n23488 ; n23489
g23234 and n7677 n8365 ; n23490
g23235 and n23489 n23490_not ; n23491
g23236 and a[50] n23491_not ; n23492
g23237 and a[50] n23492_not ; n23493
g23238 and n23491_not n23492_not ; n23494
g23239 and n23493_not n23494_not ; n23495
g23240 and n23484 n23495_not ; n23496
g23241 and n23484 n23496_not ; n23497
g23242 and n23495_not n23496_not ; n23498
g23243 and n23497_not n23498_not ; n23499
g23244 and n23261_not n23265_not ; n23500
g23245 and n23499 n23500 ; n23501
g23246 and n23499_not n23500_not ; n23502
g23247 and n23501_not n23502_not ; n23503
g23248 and b[49] n7446 ; n23504
g23249 and b[47] n7787 ; n23505
g23250 and b[48] n7441 ; n23506
g23251 and n23505_not n23506_not ; n23507
g23252 and n23504_not n23507 ; n23508
g23253 and n7449 n8625 ; n23509
g23254 and n23508 n23509_not ; n23510
g23255 and a[47] n23510_not ; n23511
g23256 and a[47] n23511_not ; n23512
g23257 and n23510_not n23511_not ; n23513
g23258 and n23512_not n23513_not ; n23514
g23259 and n23503 n23514_not ; n23515
g23260 and n23503 n23515_not ; n23516
g23261 and n23514_not n23515_not ; n23517
g23262 and n23516_not n23517_not ; n23518
g23263 and n23278_not n23284_not ; n23519
g23264 and n23518 n23519 ; n23520
g23265 and n23518_not n23519_not ; n23521
g23266 and n23520_not n23521_not ; n23522
g23267 and b[52] n6595 ; n23523
g23268 and b[50] n6902 ; n23524
g23269 and b[51] n6590 ; n23525
g23270 and n23524_not n23525_not ; n23526
g23271 and n23523_not n23526 ; n23527
g23272 and n6598 n9628 ; n23528
g23273 and n23527 n23528_not ; n23529
g23274 and a[44] n23529_not ; n23530
g23275 and a[44] n23530_not ; n23531
g23276 and n23529_not n23530_not ; n23532
g23277 and n23531_not n23532_not ; n23533
g23278 and n23522 n23533_not ; n23534
g23279 and n23522 n23534_not ; n23535
g23280 and n23533_not n23534_not ; n23536
g23281 and n23535_not n23536_not ; n23537
g23282 and n23302_not n23537 ; n23538
g23283 and n23302 n23537_not ; n23539
g23284 and n23538_not n23539_not ; n23540
g23285 and b[55] n5777 ; n23541
g23286 and b[53] n6059 ; n23542
g23287 and b[54] n5772 ; n23543
g23288 and n23542_not n23543_not ; n23544
g23289 and n23541_not n23544 ; n23545
g23290 and n5780 n10684 ; n23546
g23291 and n23545 n23546_not ; n23547
g23292 and a[41] n23547_not ; n23548
g23293 and a[41] n23548_not ; n23549
g23294 and n23547_not n23548_not ; n23550
g23295 and n23549_not n23550_not ; n23551
g23296 and n23540_not n23551_not ; n23552
g23297 and n23540 n23551 ; n23553
g23298 and n23552_not n23553_not ; n23554
g23299 and n23398_not n23554 ; n23555
g23300 and n23398 n23554_not ; n23556
g23301 and n23555_not n23556_not ; n23557
g23302 and n23397_not n23557 ; n23558
g23303 and n23557 n23558_not ; n23559
g23304 and n23397_not n23558_not ; n23560
g23305 and n23559_not n23560_not ; n23561
g23306 and n23322_not n23328_not ; n23562
g23307 and n23561 n23562 ; n23563
g23308 and n23561_not n23562_not ; n23564
g23309 and n23563_not n23564_not ; n23565
g23310 and b[61] n4287 ; n23566
g23311 and b[59] n4532 ; n23567
g23312 and b[60] n4282 ; n23568
g23313 and n23567_not n23568_not ; n23569
g23314 and n23566_not n23569 ; n23570
g23315 and n4290 n12969 ; n23571
g23316 and n23570 n23571_not ; n23572
g23317 and a[35] n23572_not ; n23573
g23318 and a[35] n23573_not ; n23574
g23319 and n23572_not n23573_not ; n23575
g23320 and n23574_not n23575_not ; n23576
g23321 and n23565 n23576_not ; n23577
g23322 and n23565_not n23576 ; n23578
g23323 and n23386 n23578_not ; n23579
g23324 and n23577_not n23579 ; n23580
g23325 and n23386 n23580_not ; n23581
g23326 and n23578_not n23580_not ; n23582
g23327 and n23577_not n23582 ; n23583
g23328 and n23581_not n23583_not ; n23584
g23329 and n23361_not n23366_not ; n23585
g23330 and n23584_not n23585_not ; n23586
g23331 and n23584_not n23586_not ; n23587
g23332 and n23585_not n23586_not ; n23588
g23333 and n23587_not n23588_not ; n23589
g23334 and n23368_not n23371_not ; n23590
g23335 and n23589_not n23590_not ; n23591
g23336 and n23589 n23590 ; n23592
g23337 and n23591_not n23592_not ; f[94]
g23338 and n23586_not n23591_not ; n23594
g23339 and n23384_not n23580_not ; n23595
g23340 and n23564_not n23577_not ; n23596
g23341 and b[63] n3843 ; n23597
g23342 and n3641 n13797 ; n23598
g23343 and n23597_not n23598_not ; n23599
g23344 and a[32] n23599_not ; n23600
g23345 and a[32] n23600_not ; n23601
g23346 and n23599_not n23600_not ; n23602
g23347 and n23601_not n23602_not ; n23603
g23348 and n23596_not n23603_not ; n23604
g23349 and n23596_not n23604_not ; n23605
g23350 and n23603_not n23604_not ; n23606
g23351 and n23605_not n23606_not ; n23607
g23352 and n23302_not n23537_not ; n23608
g23353 and n23552_not n23608_not ; n23609
g23354 and b[56] n5777 ; n23610
g23355 and b[54] n6059 ; n23611
g23356 and b[55] n5772 ; n23612
g23357 and n23611_not n23612_not ; n23613
g23358 and n23610_not n23613 ; n23614
g23359 and n5780 n10708 ; n23615
g23360 and n23614 n23615_not ; n23616
g23361 and a[41] n23616_not ; n23617
g23362 and a[41] n23617_not ; n23618
g23363 and n23616_not n23617_not ; n23619
g23364 and n23618_not n23619_not ; n23620
g23365 and n23521_not n23534_not ; n23621
g23366 and b[53] n6595 ; n23622
g23367 and b[51] n6902 ; n23623
g23368 and b[52] n6590 ; n23624
g23369 and n23623_not n23624_not ; n23625
g23370 and n23622_not n23625 ; n23626
g23371 and n6598 n9972 ; n23627
g23372 and n23626 n23627_not ; n23628
g23373 and a[44] n23628_not ; n23629
g23374 and a[44] n23629_not ; n23630
g23375 and n23628_not n23629_not ; n23631
g23376 and n23630_not n23631_not ; n23632
g23377 and n23502_not n23515_not ; n23633
g23378 and n23473_not n23476_not ; n23634
g23379 and b[44] n9339 ; n23635
g23380 and b[42] n9732 ; n23636
g23381 and b[43] n9334 ; n23637
g23382 and n23636_not n23637_not ; n23638
g23383 and n23635_not n23638 ; n23639
g23384 and n7072 n9342 ; n23640
g23385 and n23639 n23640_not ; n23641
g23386 and a[53] n23641_not ; n23642
g23387 and a[53] n23642_not ; n23643
g23388 and n23641_not n23642_not ; n23644
g23389 and n23643_not n23644_not ; n23645
g23390 and n23465_not n23469_not ; n23646
g23391 and b[41] n10426 ; n23647
g23392 and b[39] n10796 ; n23648
g23393 and b[40] n10421 ; n23649
g23394 and n23648_not n23649_not ; n23650
g23395 and n23647_not n23650 ; n23651
g23396 and n6219 n10429 ; n23652
g23397 and n23651 n23652_not ; n23653
g23398 and a[56] n23653_not ; n23654
g23399 and a[56] n23654_not ; n23655
g23400 and n23653_not n23654_not ; n23656
g23401 and n23655_not n23656_not ; n23657
g23402 and n23457_not n23461_not ; n23658
g23403 and n23441_not n23455_not ; n23659
g23404 and b[31] n13903 ; n23660
g23405 and b[32] n13488_not ; n23661
g23406 and n23660_not n23661_not ; n23662
g23407 and n23438_not n23662 ; n23663
g23408 and n23438 n23662_not ; n23664
g23409 and n23659_not n23664_not ; n23665
g23410 and n23663_not n23665 ; n23666
g23411 and n23659_not n23666_not ; n23667
g23412 and n23663_not n23666_not ; n23668
g23413 and n23664_not n23668 ; n23669
g23414 and n23667_not n23669_not ; n23670
g23415 and b[35] n12668 ; n23671
g23416 and b[33] n13047 ; n23672
g23417 and b[34] n12663 ; n23673
g23418 and n23672_not n23673_not ; n23674
g23419 and n23671_not n23674 ; n23675
g23420 and n4696 n12671 ; n23676
g23421 and n23675 n23676_not ; n23677
g23422 and a[62] n23677_not ; n23678
g23423 and a[62] n23678_not ; n23679
g23424 and n23677_not n23678_not ; n23680
g23425 and n23679_not n23680_not ; n23681
g23426 and n23670_not n23681_not ; n23682
g23427 and n23670_not n23682_not ; n23683
g23428 and n23681_not n23682_not ; n23684
g23429 and n23683_not n23684_not ; n23685
g23430 and b[38] n11531 ; n23686
g23431 and b[36] n11896 ; n23687
g23432 and b[37] n11526 ; n23688
g23433 and n23687_not n23688_not ; n23689
g23434 and n23686_not n23689 ; n23690
g23435 and n5205 n11534 ; n23691
g23436 and n23690 n23691_not ; n23692
g23437 and a[59] n23692_not ; n23693
g23438 and a[59] n23693_not ; n23694
g23439 and n23692_not n23693_not ; n23695
g23440 and n23694_not n23695_not ; n23696
g23441 and n23685_not n23696 ; n23697
g23442 and n23685 n23696_not ; n23698
g23443 and n23697_not n23698_not ; n23699
g23444 and n23658_not n23699_not ; n23700
g23445 and n23658 n23699 ; n23701
g23446 and n23700_not n23701_not ; n23702
g23447 and n23657_not n23702 ; n23703
g23448 and n23657 n23702_not ; n23704
g23449 and n23703_not n23704_not ; n23705
g23450 and n23646_not n23705 ; n23706
g23451 and n23646 n23705_not ; n23707
g23452 and n23706_not n23707_not ; n23708
g23453 and n23645_not n23708 ; n23709
g23454 and n23645 n23708_not ; n23710
g23455 and n23709_not n23710_not ; n23711
g23456 and n23634_not n23711 ; n23712
g23457 and n23634 n23711_not ; n23713
g23458 and n23712_not n23713_not ; n23714
g23459 and b[47] n8362 ; n23715
g23460 and b[45] n8715 ; n23716
g23461 and b[46] n8357 ; n23717
g23462 and n23716_not n23717_not ; n23718
g23463 and n23715_not n23718 ; n23719
g23464 and n7703 n8365 ; n23720
g23465 and n23719 n23720_not ; n23721
g23466 and a[50] n23721_not ; n23722
g23467 and a[50] n23722_not ; n23723
g23468 and n23721_not n23722_not ; n23724
g23469 and n23723_not n23724_not ; n23725
g23470 and n23714 n23725_not ; n23726
g23471 and n23714 n23726_not ; n23727
g23472 and n23725_not n23726_not ; n23728
g23473 and n23727_not n23728_not ; n23729
g23474 and n23483_not n23496_not ; n23730
g23475 and n23729 n23730 ; n23731
g23476 and n23729_not n23730_not ; n23732
g23477 and n23731_not n23732_not ; n23733
g23478 and b[50] n7446 ; n23734
g23479 and b[48] n7787 ; n23735
g23480 and b[49] n7441 ; n23736
g23481 and n23735_not n23736_not ; n23737
g23482 and n23734_not n23737 ; n23738
g23483 and n7449 n8949 ; n23739
g23484 and n23738 n23739_not ; n23740
g23485 and a[47] n23740_not ; n23741
g23486 and a[47] n23741_not ; n23742
g23487 and n23740_not n23741_not ; n23743
g23488 and n23742_not n23743_not ; n23744
g23489 and n23733_not n23744 ; n23745
g23490 and n23733 n23744_not ; n23746
g23491 and n23745_not n23746_not ; n23747
g23492 and n23633_not n23747 ; n23748
g23493 and n23633_not n23748_not ; n23749
g23494 and n23747 n23748_not ; n23750
g23495 and n23749_not n23750_not ; n23751
g23496 and n23632_not n23751_not ; n23752
g23497 and n23632 n23750_not ; n23753
g23498 and n23749_not n23753 ; n23754
g23499 and n23752_not n23754_not ; n23755
g23500 and n23621_not n23755 ; n23756
g23501 and n23621 n23755_not ; n23757
g23502 and n23756_not n23757_not ; n23758
g23503 and n23620_not n23758 ; n23759
g23504 and n23620 n23758_not ; n23760
g23505 and n23759_not n23760_not ; n23761
g23506 and n23609_not n23761 ; n23762
g23507 and n23609 n23761_not ; n23763
g23508 and n23762_not n23763_not ; n23764
g23509 and b[59] n5035 ; n23765
g23510 and b[57] n5277 ; n23766
g23511 and b[58] n5030 ; n23767
g23512 and n23766_not n23767_not ; n23768
g23513 and n23765_not n23768 ; n23769
g23514 and n5038 n12179 ; n23770
g23515 and n23769 n23770_not ; n23771
g23516 and a[38] n23771_not ; n23772
g23517 and a[38] n23772_not ; n23773
g23518 and n23771_not n23772_not ; n23774
g23519 and n23773_not n23774_not ; n23775
g23520 and n23764 n23775_not ; n23776
g23521 and n23764 n23776_not ; n23777
g23522 and n23775_not n23776_not ; n23778
g23523 and n23777_not n23778_not ; n23779
g23524 and n23555_not n23558_not ; n23780
g23525 and n23779 n23780 ; n23781
g23526 and n23779_not n23780_not ; n23782
g23527 and n23781_not n23782_not ; n23783
g23528 and b[62] n4287 ; n23784
g23529 and b[60] n4532 ; n23785
g23530 and b[61] n4282 ; n23786
g23531 and n23785_not n23786_not ; n23787
g23532 and n23784_not n23787 ; n23788
g23533 and n4290 n13370 ; n23789
g23534 and n23788 n23789_not ; n23790
g23535 and a[35] n23790_not ; n23791
g23536 and a[35] n23791_not ; n23792
g23537 and n23790_not n23791_not ; n23793
g23538 and n23792_not n23793_not ; n23794
g23539 and n23783 n23794_not ; n23795
g23540 and n23783 n23795_not ; n23796
g23541 and n23794_not n23795_not ; n23797
g23542 and n23796_not n23797_not ; n23798
g23543 and n23607_not n23798 ; n23799
g23544 and n23607 n23798_not ; n23800
g23545 and n23799_not n23800_not ; n23801
g23546 and n23595_not n23801_not ; n23802
g23547 and n23595_not n23802_not ; n23803
g23548 and n23801_not n23802_not ; n23804
g23549 and n23803_not n23804_not ; n23805
g23550 and n23594_not n23805_not ; n23806
g23551 and n23594 n23804_not ; n23807
g23552 and n23803_not n23807 ; n23808
g23553 and n23806_not n23808_not ; f[95]
g23554 and n23802_not n23806_not ; n23810
g23555 and n23607_not n23798_not ; n23811
g23556 and n23604_not n23811_not ; n23812
g23557 and b[57] n5777 ; n23813
g23558 and b[55] n6059 ; n23814
g23559 and b[56] n5772 ; n23815
g23560 and n23814_not n23815_not ; n23816
g23561 and n23813_not n23816 ; n23817
g23562 and n5780 n11410 ; n23818
g23563 and n23817 n23818_not ; n23819
g23564 and a[41] n23819_not ; n23820
g23565 and a[41] n23820_not ; n23821
g23566 and n23819_not n23820_not ; n23822
g23567 and n23821_not n23822_not ; n23823
g23568 and n23748_not n23752_not ; n23824
g23569 and n23732_not n23746_not ; n23825
g23570 and b[42] n10426 ; n23826
g23571 and b[40] n10796 ; n23827
g23572 and b[41] n10421 ; n23828
g23573 and n23827_not n23828_not ; n23829
g23574 and n23826_not n23829 ; n23830
g23575 and n6489 n10429 ; n23831
g23576 and n23830 n23831_not ; n23832
g23577 and a[56] n23832_not ; n23833
g23578 and a[56] n23833_not ; n23834
g23579 and n23832_not n23833_not ; n23835
g23580 and n23834_not n23835_not ; n23836
g23581 and n23685_not n23696_not ; n23837
g23582 and n23682_not n23837_not ; n23838
g23583 and b[32] n13903 ; n23839
g23584 and b[33] n13488_not ; n23840
g23585 and n23839_not n23840_not ; n23841
g23586 and a[32]_not n23841_not ; n23842
g23587 and a[32] n23841 ; n23843
g23588 and n23842_not n23843_not ; n23844
g23589 and n23662_not n23844 ; n23845
g23590 and n23662_not n23845_not ; n23846
g23591 and n23844 n23845_not ; n23847
g23592 and n23846_not n23847_not ; n23848
g23593 and n23668_not n23848_not ; n23849
g23594 and n23668_not n23849_not ; n23850
g23595 and n23848_not n23849_not ; n23851
g23596 and n23850_not n23851_not ; n23852
g23597 and b[36] n12668 ; n23853
g23598 and b[34] n13047 ; n23854
g23599 and b[35] n12663 ; n23855
g23600 and n23854_not n23855_not ; n23856
g23601 and n23853_not n23856 ; n23857
g23602 and n4922 n12671 ; n23858
g23603 and n23857 n23858_not ; n23859
g23604 and a[62] n23859_not ; n23860
g23605 and a[62] n23860_not ; n23861
g23606 and n23859_not n23860_not ; n23862
g23607 and n23861_not n23862_not ; n23863
g23608 and n23852_not n23863 ; n23864
g23609 and n23852 n23863_not ; n23865
g23610 and n23864_not n23865_not ; n23866
g23611 and b[39] n11531 ; n23867
g23612 and b[37] n11896 ; n23868
g23613 and b[38] n11526 ; n23869
g23614 and n23868_not n23869_not ; n23870
g23615 and n23867_not n23870 ; n23871
g23616 and n5451 n11534 ; n23872
g23617 and n23871 n23872_not ; n23873
g23618 and a[59] n23873_not ; n23874
g23619 and a[59] n23874_not ; n23875
g23620 and n23873_not n23874_not ; n23876
g23621 and n23875_not n23876_not ; n23877
g23622 and n23866_not n23877_not ; n23878
g23623 and n23866 n23877 ; n23879
g23624 and n23878_not n23879_not ; n23880
g23625 and n23838_not n23880 ; n23881
g23626 and n23838 n23880_not ; n23882
g23627 and n23881_not n23882_not ; n23883
g23628 and n23836_not n23883 ; n23884
g23629 and n23883 n23884_not ; n23885
g23630 and n23836_not n23884_not ; n23886
g23631 and n23885_not n23886_not ; n23887
g23632 and n23700_not n23703_not ; n23888
g23633 and n23887 n23888 ; n23889
g23634 and n23887_not n23888_not ; n23890
g23635 and n23889_not n23890_not ; n23891
g23636 and b[45] n9339 ; n23892
g23637 and b[43] n9732 ; n23893
g23638 and b[44] n9334 ; n23894
g23639 and n23893_not n23894_not ; n23895
g23640 and n23892_not n23895 ; n23896
g23641 and n7361 n9342 ; n23897
g23642 and n23896 n23897_not ; n23898
g23643 and a[53] n23898_not ; n23899
g23644 and a[53] n23899_not ; n23900
g23645 and n23898_not n23899_not ; n23901
g23646 and n23900_not n23901_not ; n23902
g23647 and n23891 n23902_not ; n23903
g23648 and n23891 n23903_not ; n23904
g23649 and n23902_not n23903_not ; n23905
g23650 and n23904_not n23905_not ; n23906
g23651 and n23706_not n23709_not ; n23907
g23652 and n23906 n23907 ; n23908
g23653 and n23906_not n23907_not ; n23909
g23654 and n23908_not n23909_not ; n23910
g23655 and b[48] n8362 ; n23911
g23656 and b[46] n8715 ; n23912
g23657 and b[47] n8357 ; n23913
g23658 and n23912_not n23913_not ; n23914
g23659 and n23911_not n23914 ; n23915
g23660 and n8009 n8365 ; n23916
g23661 and n23915 n23916_not ; n23917
g23662 and a[50] n23917_not ; n23918
g23663 and a[50] n23918_not ; n23919
g23664 and n23917_not n23918_not ; n23920
g23665 and n23919_not n23920_not ; n23921
g23666 and n23910 n23921_not ; n23922
g23667 and n23910 n23922_not ; n23923
g23668 and n23921_not n23922_not ; n23924
g23669 and n23923_not n23924_not ; n23925
g23670 and n23712_not n23726_not ; n23926
g23671 and n23925 n23926 ; n23927
g23672 and n23925_not n23926_not ; n23928
g23673 and n23927_not n23928_not ; n23929
g23674 and b[51] n7446 ; n23930
g23675 and b[49] n7787 ; n23931
g23676 and b[50] n7441 ; n23932
g23677 and n23931_not n23932_not ; n23933
g23678 and n23930_not n23933 ; n23934
g23679 and n7449 n8976 ; n23935
g23680 and n23934 n23935_not ; n23936
g23681 and a[47] n23936_not ; n23937
g23682 and a[47] n23937_not ; n23938
g23683 and n23936_not n23937_not ; n23939
g23684 and n23938_not n23939_not ; n23940
g23685 and n23929 n23940_not ; n23941
g23686 and n23929_not n23940 ; n23942
g23687 and n23825_not n23942_not ; n23943
g23688 and n23941_not n23943 ; n23944
g23689 and n23825_not n23944_not ; n23945
g23690 and n23941_not n23944_not ; n23946
g23691 and n23942_not n23946 ; n23947
g23692 and n23945_not n23947_not ; n23948
g23693 and b[54] n6595 ; n23949
g23694 and b[52] n6902 ; n23950
g23695 and b[53] n6590 ; n23951
g23696 and n23950_not n23951_not ; n23952
g23697 and n23949_not n23952 ; n23953
g23698 and n6598 n9998 ; n23954
g23699 and n23953 n23954_not ; n23955
g23700 and a[44] n23955_not ; n23956
g23701 and a[44] n23956_not ; n23957
g23702 and n23955_not n23956_not ; n23958
g23703 and n23957_not n23958_not ; n23959
g23704 and n23948 n23959 ; n23960
g23705 and n23948_not n23959_not ; n23961
g23706 and n23960_not n23961_not ; n23962
g23707 and n23824_not n23962 ; n23963
g23708 and n23824 n23962_not ; n23964
g23709 and n23963_not n23964_not ; n23965
g23710 and n23823_not n23965 ; n23966
g23711 and n23965 n23966_not ; n23967
g23712 and n23823_not n23966_not ; n23968
g23713 and n23967_not n23968_not ; n23969
g23714 and n23756_not n23759_not ; n23970
g23715 and n23969 n23970 ; n23971
g23716 and n23969_not n23970_not ; n23972
g23717 and n23971_not n23972_not ; n23973
g23718 and b[60] n5035 ; n23974
g23719 and b[58] n5277 ; n23975
g23720 and b[59] n5030 ; n23976
g23721 and n23975_not n23976_not ; n23977
g23722 and n23974_not n23977 ; n23978
g23723 and n5038 n12211 ; n23979
g23724 and n23978 n23979_not ; n23980
g23725 and a[38] n23980_not ; n23981
g23726 and a[38] n23981_not ; n23982
g23727 and n23980_not n23981_not ; n23983
g23728 and n23982_not n23983_not ; n23984
g23729 and n23973 n23984_not ; n23985
g23730 and n23973 n23985_not ; n23986
g23731 and n23984_not n23985_not ; n23987
g23732 and n23986_not n23987_not ; n23988
g23733 and n23762_not n23776_not ; n23989
g23734 and n23988 n23989 ; n23990
g23735 and n23988_not n23989_not ; n23991
g23736 and n23990_not n23991_not ; n23992
g23737 and n23782_not n23795_not ; n23993
g23738 and b[63] n4287 ; n23994
g23739 and b[61] n4532 ; n23995
g23740 and b[62] n4282 ; n23996
g23741 and n23995_not n23996_not ; n23997
g23742 and n23994_not n23997 ; n23998
g23743 and n4290 n13771 ; n23999
g23744 and n23998 n23999_not ; n24000
g23745 and a[35] n24000_not ; n24001
g23746 and a[35] n24001_not ; n24002
g23747 and n24000_not n24001_not ; n24003
g23748 and n24002_not n24003_not ; n24004
g23749 and n23993_not n24004_not ; n24005
g23750 and n23993_not n24005_not ; n24006
g23751 and n24004_not n24005_not ; n24007
g23752 and n24006_not n24007_not ; n24008
g23753 and n23992_not n24008 ; n24009
g23754 and n23992 n24008_not ; n24010
g23755 and n24009_not n24010_not ; n24011
g23756 and n23812_not n24011 ; n24012
g23757 and n23812 n24011_not ; n24013
g23758 and n24012_not n24013_not ; n24014
g23759 and n23810_not n24014 ; n24015
g23760 and n23810 n24014_not ; n24016
g23761 and n24015_not n24016_not ; f[96]
g23762 and n23985_not n23991_not ; n24018
g23763 and b[62] n4532 ; n24019
g23764 and b[63] n4282 ; n24020
g23765 and n24019_not n24020_not ; n24021
g23766 and n4290_not n24021 ; n24022
g23767 and n13800 n24021 ; n24023
g23768 and n24022_not n24023_not ; n24024
g23769 and a[35] n24024_not ; n24025
g23770 and a[35]_not n24024 ; n24026
g23771 and n24025_not n24026_not ; n24027
g23772 and n24018_not n24027_not ; n24028
g23773 and n24018 n24027 ; n24029
g23774 and n24028_not n24029_not ; n24030
g23775 and b[58] n5777 ; n24031
g23776 and b[56] n6059 ; n24032
g23777 and b[57] n5772 ; n24033
g23778 and n24032_not n24033_not ; n24034
g23779 and n24031_not n24034 ; n24035
g23780 and n5780 n11436 ; n24036
g23781 and n24035 n24036_not ; n24037
g23782 and a[41] n24037_not ; n24038
g23783 and a[41] n24038_not ; n24039
g23784 and n24037_not n24038_not ; n24040
g23785 and n24039_not n24040_not ; n24041
g23786 and n23961_not n23963_not ; n24042
g23787 and b[43] n10426 ; n24043
g23788 and b[41] n10796 ; n24044
g23789 and b[42] n10421 ; n24045
g23790 and n24044_not n24045_not ; n24046
g23791 and n24043_not n24046 ; n24047
g23792 and n6515 n10429 ; n24048
g23793 and n24047 n24048_not ; n24049
g23794 and a[56] n24049_not ; n24050
g23795 and a[56] n24050_not ; n24051
g23796 and n24049_not n24050_not ; n24052
g23797 and n24051_not n24052_not ; n24053
g23798 and n23878_not n23881_not ; n24054
g23799 and b[40] n11531 ; n24055
g23800 and b[38] n11896 ; n24056
g23801 and b[39] n11526 ; n24057
g23802 and n24056_not n24057_not ; n24058
g23803 and n24055_not n24058 ; n24059
g23804 and n5955 n11534 ; n24060
g23805 and n24059 n24060_not ; n24061
g23806 and a[59] n24061_not ; n24062
g23807 and a[59] n24062_not ; n24063
g23808 and n24061_not n24062_not ; n24064
g23809 and n24063_not n24064_not ; n24065
g23810 and n23852_not n23863_not ; n24066
g23811 and n23849_not n24066_not ; n24067
g23812 and b[33] n13903 ; n24068
g23813 and b[34] n13488_not ; n24069
g23814 and n24068_not n24069_not ; n24070
g23815 and n23842_not n23845_not ; n24071
g23816 and n24070_not n24071 ; n24072
g23817 and n24070 n24071_not ; n24073
g23818 and n24072_not n24073_not ; n24074
g23819 and b[37] n12668 ; n24075
g23820 and b[35] n13047 ; n24076
g23821 and b[36] n12663 ; n24077
g23822 and n24076_not n24077_not ; n24078
g23823 and n24075_not n24078 ; n24079
g23824 and n5181 n12671 ; n24080
g23825 and n24079 n24080_not ; n24081
g23826 and a[62] n24081_not ; n24082
g23827 and a[62] n24082_not ; n24083
g23828 and n24081_not n24082_not ; n24084
g23829 and n24083_not n24084_not ; n24085
g23830 and n24074_not n24085 ; n24086
g23831 and n24074 n24085_not ; n24087
g23832 and n24086_not n24087_not ; n24088
g23833 and n24067_not n24088 ; n24089
g23834 and n24067_not n24089_not ; n24090
g23835 and n24088 n24089_not ; n24091
g23836 and n24090_not n24091_not ; n24092
g23837 and n24065_not n24092_not ; n24093
g23838 and n24065 n24091_not ; n24094
g23839 and n24090_not n24094 ; n24095
g23840 and n24093_not n24095_not ; n24096
g23841 and n24054_not n24096 ; n24097
g23842 and n24054 n24096_not ; n24098
g23843 and n24097_not n24098_not ; n24099
g23844 and n24053_not n24099 ; n24100
g23845 and n24099 n24100_not ; n24101
g23846 and n24053_not n24100_not ; n24102
g23847 and n24101_not n24102_not ; n24103
g23848 and n23884_not n23890_not ; n24104
g23849 and n24103 n24104 ; n24105
g23850 and n24103_not n24104_not ; n24106
g23851 and n24105_not n24106_not ; n24107
g23852 and b[46] n9339 ; n24108
g23853 and b[44] n9732 ; n24109
g23854 and b[45] n9334 ; n24110
g23855 and n24109_not n24110_not ; n24111
g23856 and n24108_not n24111 ; n24112
g23857 and n7677 n9342 ; n24113
g23858 and n24112 n24113_not ; n24114
g23859 and a[53] n24114_not ; n24115
g23860 and a[53] n24115_not ; n24116
g23861 and n24114_not n24115_not ; n24117
g23862 and n24116_not n24117_not ; n24118
g23863 and n24107 n24118_not ; n24119
g23864 and n24107 n24119_not ; n24120
g23865 and n24118_not n24119_not ; n24121
g23866 and n24120_not n24121_not ; n24122
g23867 and n23903_not n23909_not ; n24123
g23868 and n24122 n24123 ; n24124
g23869 and n24122_not n24123_not ; n24125
g23870 and n24124_not n24125_not ; n24126
g23871 and b[49] n8362 ; n24127
g23872 and b[47] n8715 ; n24128
g23873 and b[48] n8357 ; n24129
g23874 and n24128_not n24129_not ; n24130
g23875 and n24127_not n24130 ; n24131
g23876 and n8365 n8625 ; n24132
g23877 and n24131 n24132_not ; n24133
g23878 and a[50] n24133_not ; n24134
g23879 and a[50] n24134_not ; n24135
g23880 and n24133_not n24134_not ; n24136
g23881 and n24135_not n24136_not ; n24137
g23882 and n24126 n24137_not ; n24138
g23883 and n24126 n24138_not ; n24139
g23884 and n24137_not n24138_not ; n24140
g23885 and n24139_not n24140_not ; n24141
g23886 and n23922_not n23928_not ; n24142
g23887 and n24141 n24142 ; n24143
g23888 and n24141_not n24142_not ; n24144
g23889 and n24143_not n24144_not ; n24145
g23890 and b[52] n7446 ; n24146
g23891 and b[50] n7787 ; n24147
g23892 and b[51] n7441 ; n24148
g23893 and n24147_not n24148_not ; n24149
g23894 and n24146_not n24149 ; n24150
g23895 and n7449 n9628 ; n24151
g23896 and n24150 n24151_not ; n24152
g23897 and a[47] n24152_not ; n24153
g23898 and a[47] n24153_not ; n24154
g23899 and n24152_not n24153_not ; n24155
g23900 and n24154_not n24155_not ; n24156
g23901 and n24145 n24156_not ; n24157
g23902 and n24145 n24157_not ; n24158
g23903 and n24156_not n24157_not ; n24159
g23904 and n24158_not n24159_not ; n24160
g23905 and n23946_not n24160 ; n24161
g23906 and n23946 n24160_not ; n24162
g23907 and n24161_not n24162_not ; n24163
g23908 and b[55] n6595 ; n24164
g23909 and b[53] n6902 ; n24165
g23910 and b[54] n6590 ; n24166
g23911 and n24165_not n24166_not ; n24167
g23912 and n24164_not n24167 ; n24168
g23913 and n6598 n10684 ; n24169
g23914 and n24168 n24169_not ; n24170
g23915 and a[44] n24170_not ; n24171
g23916 and a[44] n24171_not ; n24172
g23917 and n24170_not n24171_not ; n24173
g23918 and n24172_not n24173_not ; n24174
g23919 and n24163_not n24174_not ; n24175
g23920 and n24163 n24174 ; n24176
g23921 and n24175_not n24176_not ; n24177
g23922 and n24042_not n24177 ; n24178
g23923 and n24042 n24177_not ; n24179
g23924 and n24178_not n24179_not ; n24180
g23925 and n24041_not n24180 ; n24181
g23926 and n24180 n24181_not ; n24182
g23927 and n24041_not n24181_not ; n24183
g23928 and n24182_not n24183_not ; n24184
g23929 and n23966_not n23972_not ; n24185
g23930 and n24184 n24185 ; n24186
g23931 and n24184_not n24185_not ; n24187
g23932 and n24186_not n24187_not ; n24188
g23933 and b[61] n5035 ; n24189
g23934 and b[59] n5277 ; n24190
g23935 and b[60] n5030 ; n24191
g23936 and n24190_not n24191_not ; n24192
g23937 and n24189_not n24192 ; n24193
g23938 and n5038 n12969 ; n24194
g23939 and n24193 n24194_not ; n24195
g23940 and a[38] n24195_not ; n24196
g23941 and a[38] n24196_not ; n24197
g23942 and n24195_not n24196_not ; n24198
g23943 and n24197_not n24198_not ; n24199
g23944 and n24188 n24199_not ; n24200
g23945 and n24188_not n24199 ; n24201
g23946 and n24030 n24201_not ; n24202
g23947 and n24200_not n24202 ; n24203
g23948 and n24030 n24203_not ; n24204
g23949 and n24201_not n24203_not ; n24205
g23950 and n24200_not n24205 ; n24206
g23951 and n24204_not n24206_not ; n24207
g23952 and n24005_not n24010_not ; n24208
g23953 and n24207_not n24208_not ; n24209
g23954 and n24207_not n24209_not ; n24210
g23955 and n24208_not n24209_not ; n24211
g23956 and n24210_not n24211_not ; n24212
g23957 and n24012_not n24015_not ; n24213
g23958 and n24212_not n24213_not ; n24214
g23959 and n24212 n24213 ; n24215
g23960 and n24214_not n24215_not ; f[97]
g23961 and n24209_not n24214_not ; n24217
g23962 and n24028_not n24203_not ; n24218
g23963 and n24187_not n24200_not ; n24219
g23964 and b[63] n4532 ; n24220
g23965 and n4290 n13797 ; n24221
g23966 and n24220_not n24221_not ; n24222
g23967 and a[35] n24222_not ; n24223
g23968 and a[35] n24223_not ; n24224
g23969 and n24222_not n24223_not ; n24225
g23970 and n24224_not n24225_not ; n24226
g23971 and n24219_not n24226_not ; n24227
g23972 and n24219_not n24227_not ; n24228
g23973 and n24226_not n24227_not ; n24229
g23974 and n24228_not n24229_not ; n24230
g23975 and n23946_not n24160_not ; n24231
g23976 and n24175_not n24231_not ; n24232
g23977 and b[56] n6595 ; n24233
g23978 and b[54] n6902 ; n24234
g23979 and b[55] n6590 ; n24235
g23980 and n24234_not n24235_not ; n24236
g23981 and n24233_not n24236 ; n24237
g23982 and n6598 n10708 ; n24238
g23983 and n24237 n24238_not ; n24239
g23984 and a[44] n24239_not ; n24240
g23985 and a[44] n24240_not ; n24241
g23986 and n24239_not n24240_not ; n24242
g23987 and n24241_not n24242_not ; n24243
g23988 and n24144_not n24157_not ; n24244
g23989 and b[53] n7446 ; n24245
g23990 and b[51] n7787 ; n24246
g23991 and b[52] n7441 ; n24247
g23992 and n24246_not n24247_not ; n24248
g23993 and n24245_not n24248 ; n24249
g23994 and n7449 n9972 ; n24250
g23995 and n24249 n24250_not ; n24251
g23996 and a[47] n24251_not ; n24252
g23997 and a[47] n24252_not ; n24253
g23998 and n24251_not n24252_not ; n24254
g23999 and n24253_not n24254_not ; n24255
g24000 and n24125_not n24138_not ; n24256
g24001 and n24097_not n24100_not ; n24257
g24002 and b[44] n10426 ; n24258
g24003 and b[42] n10796 ; n24259
g24004 and b[43] n10421 ; n24260
g24005 and n24259_not n24260_not ; n24261
g24006 and n24258_not n24261 ; n24262
g24007 and n7072 n10429 ; n24263
g24008 and n24262 n24263_not ; n24264
g24009 and a[56] n24264_not ; n24265
g24010 and a[56] n24265_not ; n24266
g24011 and n24264_not n24265_not ; n24267
g24012 and n24266_not n24267_not ; n24268
g24013 and n24089_not n24093_not ; n24269
g24014 and n24073_not n24087_not ; n24270
g24015 and b[34] n13903 ; n24271
g24016 and b[35] n13488_not ; n24272
g24017 and n24271_not n24272_not ; n24273
g24018 and n24070_not n24273 ; n24274
g24019 and n24070 n24273_not ; n24275
g24020 and n24270_not n24275_not ; n24276
g24021 and n24274_not n24276 ; n24277
g24022 and n24270_not n24277_not ; n24278
g24023 and n24274_not n24277_not ; n24279
g24024 and n24275_not n24279 ; n24280
g24025 and n24278_not n24280_not ; n24281
g24026 and b[38] n12668 ; n24282
g24027 and b[36] n13047 ; n24283
g24028 and b[37] n12663 ; n24284
g24029 and n24283_not n24284_not ; n24285
g24030 and n24282_not n24285 ; n24286
g24031 and n5205 n12671 ; n24287
g24032 and n24286 n24287_not ; n24288
g24033 and a[62] n24288_not ; n24289
g24034 and a[62] n24289_not ; n24290
g24035 and n24288_not n24289_not ; n24291
g24036 and n24290_not n24291_not ; n24292
g24037 and n24281_not n24292_not ; n24293
g24038 and n24281_not n24293_not ; n24294
g24039 and n24292_not n24293_not ; n24295
g24040 and n24294_not n24295_not ; n24296
g24041 and b[41] n11531 ; n24297
g24042 and b[39] n11896 ; n24298
g24043 and b[40] n11526 ; n24299
g24044 and n24298_not n24299_not ; n24300
g24045 and n24297_not n24300 ; n24301
g24046 and n6219 n11534 ; n24302
g24047 and n24301 n24302_not ; n24303
g24048 and a[59] n24303_not ; n24304
g24049 and a[59] n24304_not ; n24305
g24050 and n24303_not n24304_not ; n24306
g24051 and n24305_not n24306_not ; n24307
g24052 and n24296_not n24307 ; n24308
g24053 and n24296 n24307_not ; n24309
g24054 and n24308_not n24309_not ; n24310
g24055 and n24269_not n24310_not ; n24311
g24056 and n24269 n24310 ; n24312
g24057 and n24311_not n24312_not ; n24313
g24058 and n24268_not n24313 ; n24314
g24059 and n24268 n24313_not ; n24315
g24060 and n24314_not n24315_not ; n24316
g24061 and n24257_not n24316 ; n24317
g24062 and n24257 n24316_not ; n24318
g24063 and n24317_not n24318_not ; n24319
g24064 and b[47] n9339 ; n24320
g24065 and b[45] n9732 ; n24321
g24066 and b[46] n9334 ; n24322
g24067 and n24321_not n24322_not ; n24323
g24068 and n24320_not n24323 ; n24324
g24069 and n7703 n9342 ; n24325
g24070 and n24324 n24325_not ; n24326
g24071 and a[53] n24326_not ; n24327
g24072 and a[53] n24327_not ; n24328
g24073 and n24326_not n24327_not ; n24329
g24074 and n24328_not n24329_not ; n24330
g24075 and n24319 n24330_not ; n24331
g24076 and n24319 n24331_not ; n24332
g24077 and n24330_not n24331_not ; n24333
g24078 and n24332_not n24333_not ; n24334
g24079 and n24106_not n24119_not ; n24335
g24080 and n24334 n24335 ; n24336
g24081 and n24334_not n24335_not ; n24337
g24082 and n24336_not n24337_not ; n24338
g24083 and b[50] n8362 ; n24339
g24084 and b[48] n8715 ; n24340
g24085 and b[49] n8357 ; n24341
g24086 and n24340_not n24341_not ; n24342
g24087 and n24339_not n24342 ; n24343
g24088 and n8365 n8949 ; n24344
g24089 and n24343 n24344_not ; n24345
g24090 and a[50] n24345_not ; n24346
g24091 and a[50] n24346_not ; n24347
g24092 and n24345_not n24346_not ; n24348
g24093 and n24347_not n24348_not ; n24349
g24094 and n24338_not n24349 ; n24350
g24095 and n24338 n24349_not ; n24351
g24096 and n24350_not n24351_not ; n24352
g24097 and n24256_not n24352 ; n24353
g24098 and n24256_not n24353_not ; n24354
g24099 and n24352 n24353_not ; n24355
g24100 and n24354_not n24355_not ; n24356
g24101 and n24255_not n24356_not ; n24357
g24102 and n24255 n24355_not ; n24358
g24103 and n24354_not n24358 ; n24359
g24104 and n24357_not n24359_not ; n24360
g24105 and n24244_not n24360 ; n24361
g24106 and n24244 n24360_not ; n24362
g24107 and n24361_not n24362_not ; n24363
g24108 and n24243_not n24363 ; n24364
g24109 and n24243 n24363_not ; n24365
g24110 and n24364_not n24365_not ; n24366
g24111 and n24232_not n24366 ; n24367
g24112 and n24232 n24366_not ; n24368
g24113 and n24367_not n24368_not ; n24369
g24114 and b[59] n5777 ; n24370
g24115 and b[57] n6059 ; n24371
g24116 and b[58] n5772 ; n24372
g24117 and n24371_not n24372_not ; n24373
g24118 and n24370_not n24373 ; n24374
g24119 and n5780 n12179 ; n24375
g24120 and n24374 n24375_not ; n24376
g24121 and a[41] n24376_not ; n24377
g24122 and a[41] n24377_not ; n24378
g24123 and n24376_not n24377_not ; n24379
g24124 and n24378_not n24379_not ; n24380
g24125 and n24369 n24380_not ; n24381
g24126 and n24369 n24381_not ; n24382
g24127 and n24380_not n24381_not ; n24383
g24128 and n24382_not n24383_not ; n24384
g24129 and n24178_not n24181_not ; n24385
g24130 and n24384 n24385 ; n24386
g24131 and n24384_not n24385_not ; n24387
g24132 and n24386_not n24387_not ; n24388
g24133 and b[62] n5035 ; n24389
g24134 and b[60] n5277 ; n24390
g24135 and b[61] n5030 ; n24391
g24136 and n24390_not n24391_not ; n24392
g24137 and n24389_not n24392 ; n24393
g24138 and n5038 n13370 ; n24394
g24139 and n24393 n24394_not ; n24395
g24140 and a[38] n24395_not ; n24396
g24141 and a[38] n24396_not ; n24397
g24142 and n24395_not n24396_not ; n24398
g24143 and n24397_not n24398_not ; n24399
g24144 and n24388 n24399_not ; n24400
g24145 and n24388 n24400_not ; n24401
g24146 and n24399_not n24400_not ; n24402
g24147 and n24401_not n24402_not ; n24403
g24148 and n24230_not n24403 ; n24404
g24149 and n24230 n24403_not ; n24405
g24150 and n24404_not n24405_not ; n24406
g24151 and n24218_not n24406_not ; n24407
g24152 and n24218 n24406 ; n24408
g24153 and n24407_not n24408_not ; n24409
g24154 and n24217_not n24409 ; n24410
g24155 and n24217 n24409_not ; n24411
g24156 and n24410_not n24411_not ; f[98]
g24157 and n24407_not n24410_not ; n24413
g24158 and n24353_not n24357_not ; n24414
g24159 and b[54] n7446 ; n24415
g24160 and b[52] n7787 ; n24416
g24161 and b[53] n7441 ; n24417
g24162 and n24416_not n24417_not ; n24418
g24163 and n24415_not n24418 ; n24419
g24164 and n7449 n9998 ; n24420
g24165 and n24419 n24420_not ; n24421
g24166 and a[47] n24421_not ; n24422
g24167 and a[47] n24422_not ; n24423
g24168 and n24421_not n24422_not ; n24424
g24169 and n24423_not n24424_not ; n24425
g24170 and n24337_not n24351_not ; n24426
g24171 and b[35] n13903 ; n24427
g24172 and b[36] n13488_not ; n24428
g24173 and n24427_not n24428_not ; n24429
g24174 and a[35] n24273_not ; n24430
g24175 and a[35]_not n24273 ; n24431
g24176 and n24430_not n24431_not ; n24432
g24177 and n24429_not n24432_not ; n24433
g24178 and n24429 n24432 ; n24434
g24179 and n24433_not n24434_not ; n24435
g24180 and n24279_not n24435 ; n24436
g24181 and n24279 n24435_not ; n24437
g24182 and n24436_not n24437_not ; n24438
g24183 and b[39] n12668 ; n24439
g24184 and b[37] n13047 ; n24440
g24185 and b[38] n12663 ; n24441
g24186 and n24440_not n24441_not ; n24442
g24187 and n24439_not n24442 ; n24443
g24188 and n5451 n12671 ; n24444
g24189 and n24443 n24444_not ; n24445
g24190 and a[62] n24445_not ; n24446
g24191 and a[62] n24446_not ; n24447
g24192 and n24445_not n24446_not ; n24448
g24193 and n24447_not n24448_not ; n24449
g24194 and n24438_not n24449 ; n24450
g24195 and n24438 n24449_not ; n24451
g24196 and n24450_not n24451_not ; n24452
g24197 and b[42] n11531 ; n24453
g24198 and b[40] n11896 ; n24454
g24199 and b[41] n11526 ; n24455
g24200 and n24454_not n24455_not ; n24456
g24201 and n24453_not n24456 ; n24457
g24202 and n6489 n11534 ; n24458
g24203 and n24457 n24458_not ; n24459
g24204 and a[59] n24459_not ; n24460
g24205 and a[59] n24460_not ; n24461
g24206 and n24459_not n24460_not ; n24462
g24207 and n24461_not n24462_not ; n24463
g24208 and n24452 n24463_not ; n24464
g24209 and n24452 n24464_not ; n24465
g24210 and n24463_not n24464_not ; n24466
g24211 and n24465_not n24466_not ; n24467
g24212 and n24296_not n24307_not ; n24468
g24213 and n24293_not n24468_not ; n24469
g24214 and n24467_not n24469_not ; n24470
g24215 and n24467_not n24470_not ; n24471
g24216 and n24469_not n24470_not ; n24472
g24217 and n24471_not n24472_not ; n24473
g24218 and b[45] n10426 ; n24474
g24219 and b[43] n10796 ; n24475
g24220 and b[44] n10421 ; n24476
g24221 and n24475_not n24476_not ; n24477
g24222 and n24474_not n24477 ; n24478
g24223 and n7361 n10429 ; n24479
g24224 and n24478 n24479_not ; n24480
g24225 and a[56] n24480_not ; n24481
g24226 and a[56] n24481_not ; n24482
g24227 and n24480_not n24481_not ; n24483
g24228 and n24482_not n24483_not ; n24484
g24229 and n24473_not n24484_not ; n24485
g24230 and n24473_not n24485_not ; n24486
g24231 and n24484_not n24485_not ; n24487
g24232 and n24486_not n24487_not ; n24488
g24233 and n24311_not n24314_not ; n24489
g24234 and n24488 n24489 ; n24490
g24235 and n24488_not n24489_not ; n24491
g24236 and n24490_not n24491_not ; n24492
g24237 and b[48] n9339 ; n24493
g24238 and b[46] n9732 ; n24494
g24239 and b[47] n9334 ; n24495
g24240 and n24494_not n24495_not ; n24496
g24241 and n24493_not n24496 ; n24497
g24242 and n8009 n9342 ; n24498
g24243 and n24497 n24498_not ; n24499
g24244 and a[53] n24499_not ; n24500
g24245 and a[53] n24500_not ; n24501
g24246 and n24499_not n24500_not ; n24502
g24247 and n24501_not n24502_not ; n24503
g24248 and n24492 n24503_not ; n24504
g24249 and n24492 n24504_not ; n24505
g24250 and n24503_not n24504_not ; n24506
g24251 and n24505_not n24506_not ; n24507
g24252 and n24317_not n24331_not ; n24508
g24253 and n24507 n24508 ; n24509
g24254 and n24507_not n24508_not ; n24510
g24255 and n24509_not n24510_not ; n24511
g24256 and b[51] n8362 ; n24512
g24257 and b[49] n8715 ; n24513
g24258 and b[50] n8357 ; n24514
g24259 and n24513_not n24514_not ; n24515
g24260 and n24512_not n24515 ; n24516
g24261 and n8365 n8976 ; n24517
g24262 and n24516 n24517_not ; n24518
g24263 and a[50] n24518_not ; n24519
g24264 and a[50] n24519_not ; n24520
g24265 and n24518_not n24519_not ; n24521
g24266 and n24520_not n24521_not ; n24522
g24267 and n24511_not n24522 ; n24523
g24268 and n24511 n24522_not ; n24524
g24269 and n24523_not n24524_not ; n24525
g24270 and n24426_not n24525 ; n24526
g24271 and n24426 n24525_not ; n24527
g24272 and n24526_not n24527_not ; n24528
g24273 and n24425_not n24528 ; n24529
g24274 and n24425 n24528_not ; n24530
g24275 and n24529_not n24530_not ; n24531
g24276 and n24414_not n24531 ; n24532
g24277 and n24414 n24531_not ; n24533
g24278 and n24532_not n24533_not ; n24534
g24279 and b[57] n6595 ; n24535
g24280 and b[55] n6902 ; n24536
g24281 and b[56] n6590 ; n24537
g24282 and n24536_not n24537_not ; n24538
g24283 and n24535_not n24538 ; n24539
g24284 and n6598 n11410 ; n24540
g24285 and n24539 n24540_not ; n24541
g24286 and a[44] n24541_not ; n24542
g24287 and a[44] n24542_not ; n24543
g24288 and n24541_not n24542_not ; n24544
g24289 and n24543_not n24544_not ; n24545
g24290 and n24534 n24545_not ; n24546
g24291 and n24534 n24546_not ; n24547
g24292 and n24545_not n24546_not ; n24548
g24293 and n24547_not n24548_not ; n24549
g24294 and n24361_not n24364_not ; n24550
g24295 and n24549 n24550 ; n24551
g24296 and n24549_not n24550_not ; n24552
g24297 and n24551_not n24552_not ; n24553
g24298 and b[60] n5777 ; n24554
g24299 and b[58] n6059 ; n24555
g24300 and b[59] n5772 ; n24556
g24301 and n24555_not n24556_not ; n24557
g24302 and n24554_not n24557 ; n24558
g24303 and n5780 n12211 ; n24559
g24304 and n24558 n24559_not ; n24560
g24305 and a[41] n24560_not ; n24561
g24306 and a[41] n24561_not ; n24562
g24307 and n24560_not n24561_not ; n24563
g24308 and n24562_not n24563_not ; n24564
g24309 and n24553 n24564_not ; n24565
g24310 and n24553 n24565_not ; n24566
g24311 and n24564_not n24565_not ; n24567
g24312 and n24566_not n24567_not ; n24568
g24313 and n24367_not n24381_not ; n24569
g24314 and n24568 n24569 ; n24570
g24315 and n24568_not n24569_not ; n24571
g24316 and n24570_not n24571_not ; n24572
g24317 and b[63] n5035 ; n24573
g24318 and b[61] n5277 ; n24574
g24319 and b[62] n5030 ; n24575
g24320 and n24574_not n24575_not ; n24576
g24321 and n24573_not n24576 ; n24577
g24322 and n5038 n13771 ; n24578
g24323 and n24577 n24578_not ; n24579
g24324 and a[38] n24579_not ; n24580
g24325 and a[38] n24580_not ; n24581
g24326 and n24579_not n24580_not ; n24582
g24327 and n24581_not n24582_not ; n24583
g24328 and n24572 n24583_not ; n24584
g24329 and n24572 n24584_not ; n24585
g24330 and n24583_not n24584_not ; n24586
g24331 and n24585_not n24586_not ; n24587
g24332 and n24387_not n24400_not ; n24588
g24333 and n24587 n24588 ; n24589
g24334 and n24587_not n24588_not ; n24590
g24335 and n24589_not n24590_not ; n24591
g24336 and n24230_not n24403_not ; n24592
g24337 and n24227_not n24592_not ; n24593
g24338 and n24591 n24593_not ; n24594
g24339 and n24591_not n24593 ; n24595
g24340 and n24594_not n24595_not ; n24596
g24341 and n24413_not n24596 ; n24597
g24342 and n24413 n24596_not ; n24598
g24343 and n24597_not n24598_not ; f[99]
g24344 and n24565_not n24571_not ; n24600
g24345 and b[62] n5277 ; n24601
g24346 and b[63] n5030 ; n24602
g24347 and n24601_not n24602_not ; n24603
g24348 and n5038_not n24603 ; n24604
g24349 and n13800 n24603 ; n24605
g24350 and n24604_not n24605_not ; n24606
g24351 and a[38] n24606_not ; n24607
g24352 and a[38]_not n24606 ; n24608
g24353 and n24607_not n24608_not ; n24609
g24354 and n24600_not n24609_not ; n24610
g24355 and n24600 n24609 ; n24611
g24356 and n24610_not n24611_not ; n24612
g24357 and b[40] n12668 ; n24613
g24358 and b[38] n13047 ; n24614
g24359 and b[39] n12663 ; n24615
g24360 and n24614_not n24615_not ; n24616
g24361 and n24613_not n24616 ; n24617
g24362 and n5955 n12671 ; n24618
g24363 and n24617 n24618_not ; n24619
g24364 and a[62] n24619_not ; n24620
g24365 and a[62] n24620_not ; n24621
g24366 and n24619_not n24620_not ; n24622
g24367 and n24621_not n24622_not ; n24623
g24368 and b[36] n13903 ; n24624
g24369 and b[37] n13488_not ; n24625
g24370 and n24624_not n24625_not ; n24626
g24371 and a[35]_not n24273_not ; n24627
g24372 and n24433_not n24627_not ; n24628
g24373 and n24626 n24628_not ; n24629
g24374 and n24626 n24629_not ; n24630
g24375 and n24628_not n24629_not ; n24631
g24376 and n24630_not n24631_not ; n24632
g24377 and n24623_not n24632_not ; n24633
g24378 and n24623_not n24633_not ; n24634
g24379 and n24632_not n24633_not ; n24635
g24380 and n24634_not n24635_not ; n24636
g24381 and n24436_not n24451_not ; n24637
g24382 and n24636 n24637 ; n24638
g24383 and n24636_not n24637_not ; n24639
g24384 and n24638_not n24639_not ; n24640
g24385 and b[43] n11531 ; n24641
g24386 and b[41] n11896 ; n24642
g24387 and b[42] n11526 ; n24643
g24388 and n24642_not n24643_not ; n24644
g24389 and n24641_not n24644 ; n24645
g24390 and n6515 n11534 ; n24646
g24391 and n24645 n24646_not ; n24647
g24392 and a[59] n24647_not ; n24648
g24393 and a[59] n24648_not ; n24649
g24394 and n24647_not n24648_not ; n24650
g24395 and n24649_not n24650_not ; n24651
g24396 and n24640 n24651_not ; n24652
g24397 and n24640 n24652_not ; n24653
g24398 and n24651_not n24652_not ; n24654
g24399 and n24653_not n24654_not ; n24655
g24400 and n24464_not n24470_not ; n24656
g24401 and n24655 n24656 ; n24657
g24402 and n24655_not n24656_not ; n24658
g24403 and n24657_not n24658_not ; n24659
g24404 and b[46] n10426 ; n24660
g24405 and b[44] n10796 ; n24661
g24406 and b[45] n10421 ; n24662
g24407 and n24661_not n24662_not ; n24663
g24408 and n24660_not n24663 ; n24664
g24409 and n7677 n10429 ; n24665
g24410 and n24664 n24665_not ; n24666
g24411 and a[56] n24666_not ; n24667
g24412 and a[56] n24667_not ; n24668
g24413 and n24666_not n24667_not ; n24669
g24414 and n24668_not n24669_not ; n24670
g24415 and n24659 n24670_not ; n24671
g24416 and n24659 n24671_not ; n24672
g24417 and n24670_not n24671_not ; n24673
g24418 and n24672_not n24673_not ; n24674
g24419 and n24485_not n24491_not ; n24675
g24420 and n24674 n24675 ; n24676
g24421 and n24674_not n24675_not ; n24677
g24422 and n24676_not n24677_not ; n24678
g24423 and b[49] n9339 ; n24679
g24424 and b[47] n9732 ; n24680
g24425 and b[48] n9334 ; n24681
g24426 and n24680_not n24681_not ; n24682
g24427 and n24679_not n24682 ; n24683
g24428 and n8625 n9342 ; n24684
g24429 and n24683 n24684_not ; n24685
g24430 and a[53] n24685_not ; n24686
g24431 and a[53] n24686_not ; n24687
g24432 and n24685_not n24686_not ; n24688
g24433 and n24687_not n24688_not ; n24689
g24434 and n24678 n24689_not ; n24690
g24435 and n24678 n24690_not ; n24691
g24436 and n24689_not n24690_not ; n24692
g24437 and n24691_not n24692_not ; n24693
g24438 and n24504_not n24510_not ; n24694
g24439 and n24693 n24694 ; n24695
g24440 and n24693_not n24694_not ; n24696
g24441 and n24695_not n24696_not ; n24697
g24442 and b[52] n8362 ; n24698
g24443 and b[50] n8715 ; n24699
g24444 and b[51] n8357 ; n24700
g24445 and n24699_not n24700_not ; n24701
g24446 and n24698_not n24701 ; n24702
g24447 and n8365 n9628 ; n24703
g24448 and n24702 n24703_not ; n24704
g24449 and a[50] n24704_not ; n24705
g24450 and a[50] n24705_not ; n24706
g24451 and n24704_not n24705_not ; n24707
g24452 and n24706_not n24707_not ; n24708
g24453 and n24697 n24708_not ; n24709
g24454 and n24697 n24709_not ; n24710
g24455 and n24708_not n24709_not ; n24711
g24456 and n24710_not n24711_not ; n24712
g24457 and n24524_not n24526_not ; n24713
g24458 and n24712_not n24713_not ; n24714
g24459 and n24712_not n24714_not ; n24715
g24460 and n24713_not n24714_not ; n24716
g24461 and n24715_not n24716_not ; n24717
g24462 and b[55] n7446 ; n24718
g24463 and b[53] n7787 ; n24719
g24464 and b[54] n7441 ; n24720
g24465 and n24719_not n24720_not ; n24721
g24466 and n24718_not n24721 ; n24722
g24467 and n7449 n10684 ; n24723
g24468 and n24722 n24723_not ; n24724
g24469 and a[47] n24724_not ; n24725
g24470 and a[47] n24725_not ; n24726
g24471 and n24724_not n24725_not ; n24727
g24472 and n24726_not n24727_not ; n24728
g24473 and n24717_not n24728_not ; n24729
g24474 and n24717_not n24729_not ; n24730
g24475 and n24728_not n24729_not ; n24731
g24476 and n24730_not n24731_not ; n24732
g24477 and n24529_not n24532_not ; n24733
g24478 and n24732 n24733 ; n24734
g24479 and n24732_not n24733_not ; n24735
g24480 and n24734_not n24735_not ; n24736
g24481 and b[58] n6595 ; n24737
g24482 and b[56] n6902 ; n24738
g24483 and b[57] n6590 ; n24739
g24484 and n24738_not n24739_not ; n24740
g24485 and n24737_not n24740 ; n24741
g24486 and n6598 n11436 ; n24742
g24487 and n24741 n24742_not ; n24743
g24488 and a[44] n24743_not ; n24744
g24489 and a[44] n24744_not ; n24745
g24490 and n24743_not n24744_not ; n24746
g24491 and n24745_not n24746_not ; n24747
g24492 and n24736 n24747_not ; n24748
g24493 and n24736 n24748_not ; n24749
g24494 and n24747_not n24748_not ; n24750
g24495 and n24749_not n24750_not ; n24751
g24496 and n24546_not n24552_not ; n24752
g24497 and n24751 n24752 ; n24753
g24498 and n24751_not n24752_not ; n24754
g24499 and n24753_not n24754_not ; n24755
g24500 and b[61] n5777 ; n24756
g24501 and b[59] n6059 ; n24757
g24502 and b[60] n5772 ; n24758
g24503 and n24757_not n24758_not ; n24759
g24504 and n24756_not n24759 ; n24760
g24505 and n5780 n12969 ; n24761
g24506 and n24760 n24761_not ; n24762
g24507 and a[41] n24762_not ; n24763
g24508 and a[41] n24763_not ; n24764
g24509 and n24762_not n24763_not ; n24765
g24510 and n24764_not n24765_not ; n24766
g24511 and n24755 n24766_not ; n24767
g24512 and n24755_not n24766 ; n24768
g24513 and n24612 n24768_not ; n24769
g24514 and n24767_not n24769 ; n24770
g24515 and n24612 n24770_not ; n24771
g24516 and n24768_not n24770_not ; n24772
g24517 and n24767_not n24772 ; n24773
g24518 and n24771_not n24773_not ; n24774
g24519 and n24584_not n24590_not ; n24775
g24520 and n24774 n24775 ; n24776
g24521 and n24774_not n24775_not ; n24777
g24522 and n24776_not n24777_not ; n24778
g24523 and n24594_not n24597_not ; n24779
g24524 and n24778 n24779_not ; n24780
g24525 and n24778_not n24779 ; n24781
g24526 and n24780_not n24781_not ; f[100]
g24527 and n24777_not n24780_not ; n24783
g24528 and n24610_not n24770_not ; n24784
g24529 and n24754_not n24767_not ; n24785
g24530 and b[63] n5277 ; n24786
g24531 and n5038 n13797 ; n24787
g24532 and n24786_not n24787_not ; n24788
g24533 and a[38] n24788_not ; n24789
g24534 and a[38] n24789_not ; n24790
g24535 and n24788_not n24789_not ; n24791
g24536 and n24790_not n24791_not ; n24792
g24537 and n24785_not n24792_not ; n24793
g24538 and n24785_not n24793_not ; n24794
g24539 and n24792_not n24793_not ; n24795
g24540 and n24794_not n24795_not ; n24796
g24541 and n24714_not n24729_not ; n24797
g24542 and b[56] n7446 ; n24798
g24543 and b[54] n7787 ; n24799
g24544 and b[55] n7441 ; n24800
g24545 and n24799_not n24800_not ; n24801
g24546 and n24798_not n24801 ; n24802
g24547 and n7449 n10708 ; n24803
g24548 and n24802 n24803_not ; n24804
g24549 and a[47] n24804_not ; n24805
g24550 and a[47] n24805_not ; n24806
g24551 and n24804_not n24805_not ; n24807
g24552 and n24806_not n24807_not ; n24808
g24553 and n24696_not n24709_not ; n24809
g24554 and b[53] n8362 ; n24810
g24555 and b[51] n8715 ; n24811
g24556 and b[52] n8357 ; n24812
g24557 and n24811_not n24812_not ; n24813
g24558 and n24810_not n24813 ; n24814
g24559 and n8365 n9972 ; n24815
g24560 and n24814 n24815_not ; n24816
g24561 and a[50] n24816_not ; n24817
g24562 and a[50] n24817_not ; n24818
g24563 and n24816_not n24817_not ; n24819
g24564 and n24818_not n24819_not ; n24820
g24565 and n24677_not n24690_not ; n24821
g24566 and n24629_not n24633_not ; n24822
g24567 and b[37] n13903 ; n24823
g24568 and b[38] n13488_not ; n24824
g24569 and n24823_not n24824_not ; n24825
g24570 and n24626 n24825_not ; n24826
g24571 and n24626 n24826_not ; n24827
g24572 and n24825_not n24826_not ; n24828
g24573 and n24827_not n24828_not ; n24829
g24574 and n24822_not n24829_not ; n24830
g24575 and n24822_not n24830_not ; n24831
g24576 and n24829_not n24830_not ; n24832
g24577 and n24831_not n24832_not ; n24833
g24578 and b[41] n12668 ; n24834
g24579 and b[39] n13047 ; n24835
g24580 and b[40] n12663 ; n24836
g24581 and n24835_not n24836_not ; n24837
g24582 and n24834_not n24837 ; n24838
g24583 and n6219 n12671 ; n24839
g24584 and n24838 n24839_not ; n24840
g24585 and a[62] n24840_not ; n24841
g24586 and a[62] n24841_not ; n24842
g24587 and n24840_not n24841_not ; n24843
g24588 and n24842_not n24843_not ; n24844
g24589 and n24833_not n24844_not ; n24845
g24590 and n24833_not n24845_not ; n24846
g24591 and n24844_not n24845_not ; n24847
g24592 and n24846_not n24847_not ; n24848
g24593 and b[44] n11531 ; n24849
g24594 and b[42] n11896 ; n24850
g24595 and b[43] n11526 ; n24851
g24596 and n24850_not n24851_not ; n24852
g24597 and n24849_not n24852 ; n24853
g24598 and n7072 n11534 ; n24854
g24599 and n24853 n24854_not ; n24855
g24600 and a[59] n24855_not ; n24856
g24601 and a[59] n24856_not ; n24857
g24602 and n24855_not n24856_not ; n24858
g24603 and n24857_not n24858_not ; n24859
g24604 and n24848_not n24859 ; n24860
g24605 and n24848 n24859_not ; n24861
g24606 and n24860_not n24861_not ; n24862
g24607 and n24639_not n24652_not ; n24863
g24608 and n24862 n24863 ; n24864
g24609 and n24862_not n24863_not ; n24865
g24610 and n24864_not n24865_not ; n24866
g24611 and b[47] n10426 ; n24867
g24612 and b[45] n10796 ; n24868
g24613 and b[46] n10421 ; n24869
g24614 and n24868_not n24869_not ; n24870
g24615 and n24867_not n24870 ; n24871
g24616 and n7703 n10429 ; n24872
g24617 and n24871 n24872_not ; n24873
g24618 and a[56] n24873_not ; n24874
g24619 and a[56] n24874_not ; n24875
g24620 and n24873_not n24874_not ; n24876
g24621 and n24875_not n24876_not ; n24877
g24622 and n24866 n24877_not ; n24878
g24623 and n24866 n24878_not ; n24879
g24624 and n24877_not n24878_not ; n24880
g24625 and n24879_not n24880_not ; n24881
g24626 and n24658_not n24671_not ; n24882
g24627 and n24881 n24882 ; n24883
g24628 and n24881_not n24882_not ; n24884
g24629 and n24883_not n24884_not ; n24885
g24630 and b[50] n9339 ; n24886
g24631 and b[48] n9732 ; n24887
g24632 and b[49] n9334 ; n24888
g24633 and n24887_not n24888_not ; n24889
g24634 and n24886_not n24889 ; n24890
g24635 and n8949 n9342 ; n24891
g24636 and n24890 n24891_not ; n24892
g24637 and a[53] n24892_not ; n24893
g24638 and a[53] n24893_not ; n24894
g24639 and n24892_not n24893_not ; n24895
g24640 and n24894_not n24895_not ; n24896
g24641 and n24885_not n24896 ; n24897
g24642 and n24885 n24896_not ; n24898
g24643 and n24897_not n24898_not ; n24899
g24644 and n24821_not n24899 ; n24900
g24645 and n24821_not n24900_not ; n24901
g24646 and n24899 n24900_not ; n24902
g24647 and n24901_not n24902_not ; n24903
g24648 and n24820_not n24903_not ; n24904
g24649 and n24820 n24902_not ; n24905
g24650 and n24901_not n24905 ; n24906
g24651 and n24904_not n24906_not ; n24907
g24652 and n24809_not n24907 ; n24908
g24653 and n24809 n24907_not ; n24909
g24654 and n24908_not n24909_not ; n24910
g24655 and n24808_not n24910 ; n24911
g24656 and n24808 n24910_not ; n24912
g24657 and n24911_not n24912_not ; n24913
g24658 and n24797_not n24913 ; n24914
g24659 and n24797 n24913_not ; n24915
g24660 and n24914_not n24915_not ; n24916
g24661 and b[59] n6595 ; n24917
g24662 and b[57] n6902 ; n24918
g24663 and b[58] n6590 ; n24919
g24664 and n24918_not n24919_not ; n24920
g24665 and n24917_not n24920 ; n24921
g24666 and n6598 n12179 ; n24922
g24667 and n24921 n24922_not ; n24923
g24668 and a[44] n24923_not ; n24924
g24669 and a[44] n24924_not ; n24925
g24670 and n24923_not n24924_not ; n24926
g24671 and n24925_not n24926_not ; n24927
g24672 and n24916 n24927_not ; n24928
g24673 and n24916 n24928_not ; n24929
g24674 and n24927_not n24928_not ; n24930
g24675 and n24929_not n24930_not ; n24931
g24676 and n24735_not n24748_not ; n24932
g24677 and n24931 n24932 ; n24933
g24678 and n24931_not n24932_not ; n24934
g24679 and n24933_not n24934_not ; n24935
g24680 and b[62] n5777 ; n24936
g24681 and b[60] n6059 ; n24937
g24682 and b[61] n5772 ; n24938
g24683 and n24937_not n24938_not ; n24939
g24684 and n24936_not n24939 ; n24940
g24685 and n5780 n13370 ; n24941
g24686 and n24940 n24941_not ; n24942
g24687 and a[41] n24942_not ; n24943
g24688 and a[41] n24943_not ; n24944
g24689 and n24942_not n24943_not ; n24945
g24690 and n24944_not n24945_not ; n24946
g24691 and n24935 n24946_not ; n24947
g24692 and n24935 n24947_not ; n24948
g24693 and n24946_not n24947_not ; n24949
g24694 and n24948_not n24949_not ; n24950
g24695 and n24796_not n24950 ; n24951
g24696 and n24796 n24950_not ; n24952
g24697 and n24951_not n24952_not ; n24953
g24698 and n24784_not n24953_not ; n24954
g24699 and n24784 n24953 ; n24955
g24700 and n24954_not n24955_not ; n24956
g24701 and n24783_not n24956 ; n24957
g24702 and n24783 n24956_not ; n24958
g24703 and n24957_not n24958_not ; f[101]
g24704 and n24954_not n24957_not ; n24960
g24705 and n24900_not n24904_not ; n24961
g24706 and b[54] n8362 ; n24962
g24707 and b[52] n8715 ; n24963
g24708 and b[53] n8357 ; n24964
g24709 and n24963_not n24964_not ; n24965
g24710 and n24962_not n24965 ; n24966
g24711 and n8365 n9998 ; n24967
g24712 and n24966 n24967_not ; n24968
g24713 and a[50] n24968_not ; n24969
g24714 and a[50] n24969_not ; n24970
g24715 and n24968_not n24969_not ; n24971
g24716 and n24970_not n24971_not ; n24972
g24717 and n24884_not n24898_not ; n24973
g24718 and n24826_not n24830_not ; n24974
g24719 and b[38] n13903 ; n24975
g24720 and b[39] n13488_not ; n24976
g24721 and n24975_not n24976_not ; n24977
g24722 and a[38] n24626_not ; n24978
g24723 and a[38]_not n24626 ; n24979
g24724 and n24978_not n24979_not ; n24980
g24725 and n24977_not n24980_not ; n24981
g24726 and n24977 n24980 ; n24982
g24727 and n24981_not n24982_not ; n24983
g24728 and n24974_not n24983 ; n24984
g24729 and n24974 n24983_not ; n24985
g24730 and n24984_not n24985_not ; n24986
g24731 and b[42] n12668 ; n24987
g24732 and b[40] n13047 ; n24988
g24733 and b[41] n12663 ; n24989
g24734 and n24988_not n24989_not ; n24990
g24735 and n24987_not n24990 ; n24991
g24736 and n6489 n12671 ; n24992
g24737 and n24991 n24992_not ; n24993
g24738 and a[62] n24993_not ; n24994
g24739 and a[62] n24994_not ; n24995
g24740 and n24993_not n24994_not ; n24996
g24741 and n24995_not n24996_not ; n24997
g24742 and n24986 n24997_not ; n24998
g24743 and n24986 n24998_not ; n24999
g24744 and n24997_not n24998_not ; n25000
g24745 and n24999_not n25000_not ; n25001
g24746 and b[45] n11531 ; n25002
g24747 and b[43] n11896 ; n25003
g24748 and b[44] n11526 ; n25004
g24749 and n25003_not n25004_not ; n25005
g24750 and n25002_not n25005 ; n25006
g24751 and n7361 n11534 ; n25007
g24752 and n25006 n25007_not ; n25008
g24753 and a[59] n25008_not ; n25009
g24754 and a[59] n25009_not ; n25010
g24755 and n25008_not n25009_not ; n25011
g24756 and n25010_not n25011_not ; n25012
g24757 and n25001_not n25012_not ; n25013
g24758 and n25001_not n25013_not ; n25014
g24759 and n25012_not n25013_not ; n25015
g24760 and n25014_not n25015_not ; n25016
g24761 and n24848_not n24859_not ; n25017
g24762 and n24845_not n25017_not ; n25018
g24763 and n25016_not n25018_not ; n25019
g24764 and n25016_not n25019_not ; n25020
g24765 and n25018_not n25019_not ; n25021
g24766 and n25020_not n25021_not ; n25022
g24767 and b[48] n10426 ; n25023
g24768 and b[46] n10796 ; n25024
g24769 and b[47] n10421 ; n25025
g24770 and n25024_not n25025_not ; n25026
g24771 and n25023_not n25026 ; n25027
g24772 and n8009 n10429 ; n25028
g24773 and n25027 n25028_not ; n25029
g24774 and a[56] n25029_not ; n25030
g24775 and a[56] n25030_not ; n25031
g24776 and n25029_not n25030_not ; n25032
g24777 and n25031_not n25032_not ; n25033
g24778 and n25022_not n25033_not ; n25034
g24779 and n25022_not n25034_not ; n25035
g24780 and n25033_not n25034_not ; n25036
g24781 and n25035_not n25036_not ; n25037
g24782 and n24865_not n24878_not ; n25038
g24783 and n25037 n25038 ; n25039
g24784 and n25037_not n25038_not ; n25040
g24785 and n25039_not n25040_not ; n25041
g24786 and b[51] n9339 ; n25042
g24787 and b[49] n9732 ; n25043
g24788 and b[50] n9334 ; n25044
g24789 and n25043_not n25044_not ; n25045
g24790 and n25042_not n25045 ; n25046
g24791 and n8976 n9342 ; n25047
g24792 and n25046 n25047_not ; n25048
g24793 and a[53] n25048_not ; n25049
g24794 and a[53] n25049_not ; n25050
g24795 and n25048_not n25049_not ; n25051
g24796 and n25050_not n25051_not ; n25052
g24797 and n25041_not n25052 ; n25053
g24798 and n25041 n25052_not ; n25054
g24799 and n25053_not n25054_not ; n25055
g24800 and n24973_not n25055 ; n25056
g24801 and n24973 n25055_not ; n25057
g24802 and n25056_not n25057_not ; n25058
g24803 and n24972_not n25058 ; n25059
g24804 and n24972 n25058_not ; n25060
g24805 and n25059_not n25060_not ; n25061
g24806 and n24961_not n25061 ; n25062
g24807 and n24961 n25061_not ; n25063
g24808 and n25062_not n25063_not ; n25064
g24809 and b[57] n7446 ; n25065
g24810 and b[55] n7787 ; n25066
g24811 and b[56] n7441 ; n25067
g24812 and n25066_not n25067_not ; n25068
g24813 and n25065_not n25068 ; n25069
g24814 and n7449 n11410 ; n25070
g24815 and n25069 n25070_not ; n25071
g24816 and a[47] n25071_not ; n25072
g24817 and a[47] n25072_not ; n25073
g24818 and n25071_not n25072_not ; n25074
g24819 and n25073_not n25074_not ; n25075
g24820 and n25064 n25075_not ; n25076
g24821 and n25064 n25076_not ; n25077
g24822 and n25075_not n25076_not ; n25078
g24823 and n25077_not n25078_not ; n25079
g24824 and n24908_not n24911_not ; n25080
g24825 and n25079 n25080 ; n25081
g24826 and n25079_not n25080_not ; n25082
g24827 and n25081_not n25082_not ; n25083
g24828 and b[60] n6595 ; n25084
g24829 and b[58] n6902 ; n25085
g24830 and b[59] n6590 ; n25086
g24831 and n25085_not n25086_not ; n25087
g24832 and n25084_not n25087 ; n25088
g24833 and n6598 n12211 ; n25089
g24834 and n25088 n25089_not ; n25090
g24835 and a[44] n25090_not ; n25091
g24836 and a[44] n25091_not ; n25092
g24837 and n25090_not n25091_not ; n25093
g24838 and n25092_not n25093_not ; n25094
g24839 and n25083 n25094_not ; n25095
g24840 and n25083 n25095_not ; n25096
g24841 and n25094_not n25095_not ; n25097
g24842 and n25096_not n25097_not ; n25098
g24843 and n24914_not n24928_not ; n25099
g24844 and n25098 n25099 ; n25100
g24845 and n25098_not n25099_not ; n25101
g24846 and n25100_not n25101_not ; n25102
g24847 and b[63] n5777 ; n25103
g24848 and b[61] n6059 ; n25104
g24849 and b[62] n5772 ; n25105
g24850 and n25104_not n25105_not ; n25106
g24851 and n25103_not n25106 ; n25107
g24852 and n5780 n13771 ; n25108
g24853 and n25107 n25108_not ; n25109
g24854 and a[41] n25109_not ; n25110
g24855 and a[41] n25110_not ; n25111
g24856 and n25109_not n25110_not ; n25112
g24857 and n25111_not n25112_not ; n25113
g24858 and n25102 n25113_not ; n25114
g24859 and n25102 n25114_not ; n25115
g24860 and n25113_not n25114_not ; n25116
g24861 and n25115_not n25116_not ; n25117
g24862 and n24934_not n24947_not ; n25118
g24863 and n25117 n25118 ; n25119
g24864 and n25117_not n25118_not ; n25120
g24865 and n25119_not n25120_not ; n25121
g24866 and n24796_not n24950_not ; n25122
g24867 and n24793_not n25122_not ; n25123
g24868 and n25121 n25123_not ; n25124
g24869 and n25121_not n25123 ; n25125
g24870 and n25124_not n25125_not ; n25126
g24871 and n24960_not n25126 ; n25127
g24872 and n24960 n25126_not ; n25128
g24873 and n25127_not n25128_not ; f[102]
g24874 and n25095_not n25101_not ; n25130
g24875 and b[62] n6059 ; n25131
g24876 and b[63] n5772 ; n25132
g24877 and n25131_not n25132_not ; n25133
g24878 and n5780_not n25133 ; n25134
g24879 and n13800 n25133 ; n25135
g24880 and n25134_not n25135_not ; n25136
g24881 and a[41] n25136_not ; n25137
g24882 and a[41]_not n25136 ; n25138
g24883 and n25137_not n25138_not ; n25139
g24884 and n25130_not n25139_not ; n25140
g24885 and n25130 n25139 ; n25141
g24886 and n25140_not n25141_not ; n25142
g24887 and n24984_not n24998_not ; n25143
g24888 and b[39] n13903 ; n25144
g24889 and b[40] n13488_not ; n25145
g24890 and n25144_not n25145_not ; n25146
g24891 and a[38]_not n24626_not ; n25147
g24892 and n24981_not n25147_not ; n25148
g24893 and n25146 n25148_not ; n25149
g24894 and n25146_not n25148 ; n25150
g24895 and n25149_not n25150_not ; n25151
g24896 and b[43] n12668 ; n25152
g24897 and b[41] n13047 ; n25153
g24898 and b[42] n12663 ; n25154
g24899 and n25153_not n25154_not ; n25155
g24900 and n25152_not n25155 ; n25156
g24901 and n12671_not n25156 ; n25157
g24902 and n6515_not n25156 ; n25158
g24903 and n25157_not n25158_not ; n25159
g24904 and a[62] n25159_not ; n25160
g24905 and a[62]_not n25159 ; n25161
g24906 and n25160_not n25161_not ; n25162
g24907 and n25151 n25162_not ; n25163
g24908 and n25151_not n25162 ; n25164
g24909 and n25163_not n25164_not ; n25165
g24910 and n25143_not n25165 ; n25166
g24911 and n25143 n25165_not ; n25167
g24912 and n25166_not n25167_not ; n25168
g24913 and b[46] n11531 ; n25169
g24914 and b[44] n11896 ; n25170
g24915 and b[45] n11526 ; n25171
g24916 and n25170_not n25171_not ; n25172
g24917 and n25169_not n25172 ; n25173
g24918 and n7677 n11534 ; n25174
g24919 and n25173 n25174_not ; n25175
g24920 and a[59] n25175_not ; n25176
g24921 and a[59] n25176_not ; n25177
g24922 and n25175_not n25176_not ; n25178
g24923 and n25177_not n25178_not ; n25179
g24924 and n25168 n25179_not ; n25180
g24925 and n25168 n25180_not ; n25181
g24926 and n25179_not n25180_not ; n25182
g24927 and n25181_not n25182_not ; n25183
g24928 and n25013_not n25019_not ; n25184
g24929 and n25183 n25184 ; n25185
g24930 and n25183_not n25184_not ; n25186
g24931 and n25185_not n25186_not ; n25187
g24932 and b[49] n10426 ; n25188
g24933 and b[47] n10796 ; n25189
g24934 and b[48] n10421 ; n25190
g24935 and n25189_not n25190_not ; n25191
g24936 and n25188_not n25191 ; n25192
g24937 and n8625 n10429 ; n25193
g24938 and n25192 n25193_not ; n25194
g24939 and a[56] n25194_not ; n25195
g24940 and a[56] n25195_not ; n25196
g24941 and n25194_not n25195_not ; n25197
g24942 and n25196_not n25197_not ; n25198
g24943 and n25187 n25198_not ; n25199
g24944 and n25187 n25199_not ; n25200
g24945 and n25198_not n25199_not ; n25201
g24946 and n25200_not n25201_not ; n25202
g24947 and n25034_not n25040_not ; n25203
g24948 and n25202 n25203 ; n25204
g24949 and n25202_not n25203_not ; n25205
g24950 and n25204_not n25205_not ; n25206
g24951 and b[52] n9339 ; n25207
g24952 and b[50] n9732 ; n25208
g24953 and b[51] n9334 ; n25209
g24954 and n25208_not n25209_not ; n25210
g24955 and n25207_not n25210 ; n25211
g24956 and n9342 n9628 ; n25212
g24957 and n25211 n25212_not ; n25213
g24958 and a[53] n25213_not ; n25214
g24959 and a[53] n25214_not ; n25215
g24960 and n25213_not n25214_not ; n25216
g24961 and n25215_not n25216_not ; n25217
g24962 and n25206 n25217_not ; n25218
g24963 and n25206 n25218_not ; n25219
g24964 and n25217_not n25218_not ; n25220
g24965 and n25219_not n25220_not ; n25221
g24966 and n25054_not n25056_not ; n25222
g24967 and n25221_not n25222_not ; n25223
g24968 and n25221_not n25223_not ; n25224
g24969 and n25222_not n25223_not ; n25225
g24970 and n25224_not n25225_not ; n25226
g24971 and b[55] n8362 ; n25227
g24972 and b[53] n8715 ; n25228
g24973 and b[54] n8357 ; n25229
g24974 and n25228_not n25229_not ; n25230
g24975 and n25227_not n25230 ; n25231
g24976 and n8365 n10684 ; n25232
g24977 and n25231 n25232_not ; n25233
g24978 and a[50] n25233_not ; n25234
g24979 and a[50] n25234_not ; n25235
g24980 and n25233_not n25234_not ; n25236
g24981 and n25235_not n25236_not ; n25237
g24982 and n25226_not n25237_not ; n25238
g24983 and n25226_not n25238_not ; n25239
g24984 and n25237_not n25238_not ; n25240
g24985 and n25239_not n25240_not ; n25241
g24986 and n25059_not n25062_not ; n25242
g24987 and n25241 n25242 ; n25243
g24988 and n25241_not n25242_not ; n25244
g24989 and n25243_not n25244_not ; n25245
g24990 and b[58] n7446 ; n25246
g24991 and b[56] n7787 ; n25247
g24992 and b[57] n7441 ; n25248
g24993 and n25247_not n25248_not ; n25249
g24994 and n25246_not n25249 ; n25250
g24995 and n7449 n11436 ; n25251
g24996 and n25250 n25251_not ; n25252
g24997 and a[47] n25252_not ; n25253
g24998 and a[47] n25253_not ; n25254
g24999 and n25252_not n25253_not ; n25255
g25000 and n25254_not n25255_not ; n25256
g25001 and n25245 n25256_not ; n25257
g25002 and n25245 n25257_not ; n25258
g25003 and n25256_not n25257_not ; n25259
g25004 and n25258_not n25259_not ; n25260
g25005 and n25076_not n25082_not ; n25261
g25006 and n25260 n25261 ; n25262
g25007 and n25260_not n25261_not ; n25263
g25008 and n25262_not n25263_not ; n25264
g25009 and b[61] n6595 ; n25265
g25010 and b[59] n6902 ; n25266
g25011 and b[60] n6590 ; n25267
g25012 and n25266_not n25267_not ; n25268
g25013 and n25265_not n25268 ; n25269
g25014 and n6598 n12969 ; n25270
g25015 and n25269 n25270_not ; n25271
g25016 and a[44] n25271_not ; n25272
g25017 and a[44] n25272_not ; n25273
g25018 and n25271_not n25272_not ; n25274
g25019 and n25273_not n25274_not ; n25275
g25020 and n25264 n25275_not ; n25276
g25021 and n25264_not n25275 ; n25277
g25022 and n25142 n25277_not ; n25278
g25023 and n25276_not n25278 ; n25279
g25024 and n25142 n25279_not ; n25280
g25025 and n25277_not n25279_not ; n25281
g25026 and n25276_not n25281 ; n25282
g25027 and n25280_not n25282_not ; n25283
g25028 and n25114_not n25120_not ; n25284
g25029 and n25283 n25284 ; n25285
g25030 and n25283_not n25284_not ; n25286
g25031 and n25285_not n25286_not ; n25287
g25032 and n25124_not n25127_not ; n25288
g25033 and n25287 n25288_not ; n25289
g25034 and n25287_not n25288 ; n25290
g25035 and n25289_not n25290_not ; f[103]
g25036 and n25286_not n25289_not ; n25292
g25037 and n25140_not n25279_not ; n25293
g25038 and n25263_not n25276_not ; n25294
g25039 and b[63] n6059 ; n25295
g25040 and n5780 n13797 ; n25296
g25041 and n25295_not n25296_not ; n25297
g25042 and a[41] n25297_not ; n25298
g25043 and a[41] n25298_not ; n25299
g25044 and n25297_not n25298_not ; n25300
g25045 and n25299_not n25300_not ; n25301
g25046 and n25294_not n25301_not ; n25302
g25047 and n25294_not n25302_not ; n25303
g25048 and n25301_not n25302_not ; n25304
g25049 and n25303_not n25304_not ; n25305
g25050 and b[59] n7446 ; n25306
g25051 and b[57] n7787 ; n25307
g25052 and b[58] n7441 ; n25308
g25053 and n25307_not n25308_not ; n25309
g25054 and n25306_not n25309 ; n25310
g25055 and n7449 n12179 ; n25311
g25056 and n25310 n25311_not ; n25312
g25057 and a[47] n25312_not ; n25313
g25058 and a[47] n25313_not ; n25314
g25059 and n25312_not n25313_not ; n25315
g25060 and n25314_not n25315_not ; n25316
g25061 and n25223_not n25238_not ; n25317
g25062 and b[56] n8362 ; n25318
g25063 and b[54] n8715 ; n25319
g25064 and b[55] n8357 ; n25320
g25065 and n25319_not n25320_not ; n25321
g25066 and n25318_not n25321 ; n25322
g25067 and n8365 n10708 ; n25323
g25068 and n25322 n25323_not ; n25324
g25069 and a[50] n25324_not ; n25325
g25070 and a[50] n25325_not ; n25326
g25071 and n25324_not n25325_not ; n25327
g25072 and n25326_not n25327_not ; n25328
g25073 and n25205_not n25218_not ; n25329
g25074 and b[53] n9339 ; n25330
g25075 and b[51] n9732 ; n25331
g25076 and b[52] n9334 ; n25332
g25077 and n25331_not n25332_not ; n25333
g25078 and n25330_not n25333 ; n25334
g25079 and n9342 n9972 ; n25335
g25080 and n25334 n25335_not ; n25336
g25081 and a[53] n25336_not ; n25337
g25082 and a[53] n25337_not ; n25338
g25083 and n25336_not n25337_not ; n25339
g25084 and n25338_not n25339_not ; n25340
g25085 and n25186_not n25199_not ; n25341
g25086 and n25166_not n25180_not ; n25342
g25087 and n25149_not n25163_not ; n25343
g25088 and b[40] n13903 ; n25344
g25089 and b[41] n13488_not ; n25345
g25090 and n25344_not n25345_not ; n25346
g25091 and n25146 n25346_not ; n25347
g25092 and n25146 n25347_not ; n25348
g25093 and n25346_not n25347_not ; n25349
g25094 and n25348_not n25349_not ; n25350
g25095 and n25343_not n25350_not ; n25351
g25096 and n25343_not n25351_not ; n25352
g25097 and n25350_not n25351_not ; n25353
g25098 and n25352_not n25353_not ; n25354
g25099 and b[44] n12668 ; n25355
g25100 and b[42] n13047 ; n25356
g25101 and b[43] n12663 ; n25357
g25102 and n25356_not n25357_not ; n25358
g25103 and n25355_not n25358 ; n25359
g25104 and n7072 n12671 ; n25360
g25105 and n25359 n25360_not ; n25361
g25106 and a[62] n25361_not ; n25362
g25107 and a[62] n25362_not ; n25363
g25108 and n25361_not n25362_not ; n25364
g25109 and n25363_not n25364_not ; n25365
g25110 and n25354_not n25365 ; n25366
g25111 and n25354 n25365_not ; n25367
g25112 and n25366_not n25367_not ; n25368
g25113 and b[47] n11531 ; n25369
g25114 and b[45] n11896 ; n25370
g25115 and b[46] n11526 ; n25371
g25116 and n25370_not n25371_not ; n25372
g25117 and n25369_not n25372 ; n25373
g25118 and n7703 n11534 ; n25374
g25119 and n25373 n25374_not ; n25375
g25120 and a[59] n25375_not ; n25376
g25121 and a[59] n25376_not ; n25377
g25122 and n25375_not n25376_not ; n25378
g25123 and n25377_not n25378_not ; n25379
g25124 and n25368_not n25379_not ; n25380
g25125 and n25368 n25379 ; n25381
g25126 and n25380_not n25381_not ; n25382
g25127 and n25342 n25382_not ; n25383
g25128 and n25342_not n25382 ; n25384
g25129 and n25383_not n25384_not ; n25385
g25130 and b[50] n10426 ; n25386
g25131 and b[48] n10796 ; n25387
g25132 and b[49] n10421 ; n25388
g25133 and n25387_not n25388_not ; n25389
g25134 and n25386_not n25389 ; n25390
g25135 and n8949 n10429 ; n25391
g25136 and n25390 n25391_not ; n25392
g25137 and a[56] n25392_not ; n25393
g25138 and a[56] n25393_not ; n25394
g25139 and n25392_not n25393_not ; n25395
g25140 and n25394_not n25395_not ; n25396
g25141 and n25385_not n25396 ; n25397
g25142 and n25385 n25396_not ; n25398
g25143 and n25397_not n25398_not ; n25399
g25144 and n25341_not n25399 ; n25400
g25145 and n25341_not n25400_not ; n25401
g25146 and n25399 n25400_not ; n25402
g25147 and n25401_not n25402_not ; n25403
g25148 and n25340_not n25403_not ; n25404
g25149 and n25340 n25402_not ; n25405
g25150 and n25401_not n25405 ; n25406
g25151 and n25404_not n25406_not ; n25407
g25152 and n25329_not n25407 ; n25408
g25153 and n25329_not n25408_not ; n25409
g25154 and n25407 n25408_not ; n25410
g25155 and n25409_not n25410_not ; n25411
g25156 and n25328_not n25411_not ; n25412
g25157 and n25328 n25410_not ; n25413
g25158 and n25409_not n25413 ; n25414
g25159 and n25412_not n25414_not ; n25415
g25160 and n25317_not n25415 ; n25416
g25161 and n25317 n25415_not ; n25417
g25162 and n25416_not n25417_not ; n25418
g25163 and n25316_not n25418 ; n25419
g25164 and n25418 n25419_not ; n25420
g25165 and n25316_not n25419_not ; n25421
g25166 and n25420_not n25421_not ; n25422
g25167 and n25244_not n25257_not ; n25423
g25168 and n25422 n25423 ; n25424
g25169 and n25422_not n25423_not ; n25425
g25170 and n25424_not n25425_not ; n25426
g25171 and b[62] n6595 ; n25427
g25172 and b[60] n6902 ; n25428
g25173 and b[61] n6590 ; n25429
g25174 and n25428_not n25429_not ; n25430
g25175 and n25427_not n25430 ; n25431
g25176 and n6598 n13370 ; n25432
g25177 and n25431 n25432_not ; n25433
g25178 and a[44] n25433_not ; n25434
g25179 and a[44] n25434_not ; n25435
g25180 and n25433_not n25434_not ; n25436
g25181 and n25435_not n25436_not ; n25437
g25182 and n25426 n25437_not ; n25438
g25183 and n25426 n25438_not ; n25439
g25184 and n25437_not n25438_not ; n25440
g25185 and n25439_not n25440_not ; n25441
g25186 and n25305_not n25441 ; n25442
g25187 and n25305 n25441_not ; n25443
g25188 and n25442_not n25443_not ; n25444
g25189 and n25293_not n25444_not ; n25445
g25190 and n25293 n25444 ; n25446
g25191 and n25445_not n25446_not ; n25447
g25192 and n25292_not n25447 ; n25448
g25193 and n25292 n25447_not ; n25449
g25194 and n25448_not n25449_not ; f[104]
g25195 and n25445_not n25448_not ; n25451
g25196 and b[60] n7446 ; n25452
g25197 and b[58] n7787 ; n25453
g25198 and b[59] n7441 ; n25454
g25199 and n25453_not n25454_not ; n25455
g25200 and n25452_not n25455 ; n25456
g25201 and n7449 n12211 ; n25457
g25202 and n25456 n25457_not ; n25458
g25203 and a[47] n25458_not ; n25459
g25204 and a[47] n25459_not ; n25460
g25205 and n25458_not n25459_not ; n25461
g25206 and n25460_not n25461_not ; n25462
g25207 and n25408_not n25412_not ; n25463
g25208 and b[57] n8362 ; n25464
g25209 and b[55] n8715 ; n25465
g25210 and b[56] n8357 ; n25466
g25211 and n25465_not n25466_not ; n25467
g25212 and n25464_not n25467 ; n25468
g25213 and n8365 n11410 ; n25469
g25214 and n25468 n25469_not ; n25470
g25215 and a[50] n25470_not ; n25471
g25216 and a[50] n25471_not ; n25472
g25217 and n25470_not n25471_not ; n25473
g25218 and n25472_not n25473_not ; n25474
g25219 and n25400_not n25404_not ; n25475
g25220 and n25384_not n25398_not ; n25476
g25221 and b[51] n10426 ; n25477
g25222 and b[49] n10796 ; n25478
g25223 and b[50] n10421 ; n25479
g25224 and n25478_not n25479_not ; n25480
g25225 and n25477_not n25480 ; n25481
g25226 and n8976 n10429 ; n25482
g25227 and n25481 n25482_not ; n25483
g25228 and a[56] n25483_not ; n25484
g25229 and a[56] n25484_not ; n25485
g25230 and n25483_not n25484_not ; n25486
g25231 and n25485_not n25486_not ; n25487
g25232 and a[41] n25146_not ; n25488
g25233 and a[41]_not n25146 ; n25489
g25234 and n25488_not n25489_not ; n25490
g25235 and b[41] n13903 ; n25491
g25236 and b[42] n13488_not ; n25492
g25237 and n25491_not n25492_not ; n25493
g25238 and n25490 n25493 ; n25494
g25239 and n25490_not n25493_not ; n25495
g25240 and n25494_not n25495_not ; n25496
g25241 and b[45] n12668 ; n25497
g25242 and b[43] n13047 ; n25498
g25243 and b[44] n12663 ; n25499
g25244 and n25498_not n25499_not ; n25500
g25245 and n25497_not n25500 ; n25501
g25246 and n7361 n12671 ; n25502
g25247 and n25501 n25502_not ; n25503
g25248 and a[62] n25503_not ; n25504
g25249 and a[62] n25504_not ; n25505
g25250 and n25503_not n25504_not ; n25506
g25251 and n25505_not n25506_not ; n25507
g25252 and n25496 n25507_not ; n25508
g25253 and n25496 n25508_not ; n25509
g25254 and n25507_not n25508_not ; n25510
g25255 and n25509_not n25510_not ; n25511
g25256 and n25347_not n25351_not ; n25512
g25257 and n25511 n25512 ; n25513
g25258 and n25511_not n25512_not ; n25514
g25259 and n25513_not n25514_not ; n25515
g25260 and b[48] n11531 ; n25516
g25261 and b[46] n11896 ; n25517
g25262 and b[47] n11526 ; n25518
g25263 and n25517_not n25518_not ; n25519
g25264 and n25516_not n25519 ; n25520
g25265 and n8009 n11534 ; n25521
g25266 and n25520 n25521_not ; n25522
g25267 and a[59] n25522_not ; n25523
g25268 and a[59] n25523_not ; n25524
g25269 and n25522_not n25523_not ; n25525
g25270 and n25524_not n25525_not ; n25526
g25271 and n25515 n25526_not ; n25527
g25272 and n25515 n25527_not ; n25528
g25273 and n25526_not n25527_not ; n25529
g25274 and n25528_not n25529_not ; n25530
g25275 and n25354_not n25365_not ; n25531
g25276 and n25380_not n25531_not ; n25532
g25277 and n25530_not n25532_not ; n25533
g25278 and n25530 n25532 ; n25534
g25279 and n25533_not n25534_not ; n25535
g25280 and n25487_not n25535 ; n25536
g25281 and n25487_not n25536_not ; n25537
g25282 and n25535 n25536_not ; n25538
g25283 and n25537_not n25538_not ; n25539
g25284 and n25476_not n25539_not ; n25540
g25285 and n25476_not n25540_not ; n25541
g25286 and n25539_not n25540_not ; n25542
g25287 and n25541_not n25542_not ; n25543
g25288 and b[54] n9339 ; n25544
g25289 and b[52] n9732 ; n25545
g25290 and b[53] n9334 ; n25546
g25291 and n25545_not n25546_not ; n25547
g25292 and n25544_not n25547 ; n25548
g25293 and n9342 n9998 ; n25549
g25294 and n25548 n25549_not ; n25550
g25295 and a[53] n25550_not ; n25551
g25296 and a[53] n25551_not ; n25552
g25297 and n25550_not n25551_not ; n25553
g25298 and n25552_not n25553_not ; n25554
g25299 and n25543 n25554 ; n25555
g25300 and n25543_not n25554_not ; n25556
g25301 and n25555_not n25556_not ; n25557
g25302 and n25475_not n25557 ; n25558
g25303 and n25475 n25557_not ; n25559
g25304 and n25558_not n25559_not ; n25560
g25305 and n25474 n25560_not ; n25561
g25306 and n25474_not n25560 ; n25562
g25307 and n25561_not n25562_not ; n25563
g25308 and n25463_not n25563 ; n25564
g25309 and n25463 n25563_not ; n25565
g25310 and n25564_not n25565_not ; n25566
g25311 and n25462_not n25566 ; n25567
g25312 and n25566 n25567_not ; n25568
g25313 and n25462_not n25567_not ; n25569
g25314 and n25568_not n25569_not ; n25570
g25315 and n25416_not n25419_not ; n25571
g25316 and n25570 n25571 ; n25572
g25317 and n25570_not n25571_not ; n25573
g25318 and n25572_not n25573_not ; n25574
g25319 and b[63] n6595 ; n25575
g25320 and b[61] n6902 ; n25576
g25321 and b[62] n6590 ; n25577
g25322 and n25576_not n25577_not ; n25578
g25323 and n25575_not n25578 ; n25579
g25324 and n6598 n13771 ; n25580
g25325 and n25579 n25580_not ; n25581
g25326 and a[44] n25581_not ; n25582
g25327 and a[44] n25582_not ; n25583
g25328 and n25581_not n25582_not ; n25584
g25329 and n25583_not n25584_not ; n25585
g25330 and n25574 n25585_not ; n25586
g25331 and n25574 n25586_not ; n25587
g25332 and n25585_not n25586_not ; n25588
g25333 and n25587_not n25588_not ; n25589
g25334 and n25425_not n25438_not ; n25590
g25335 and n25589 n25590 ; n25591
g25336 and n25589_not n25590_not ; n25592
g25337 and n25591_not n25592_not ; n25593
g25338 and n25305_not n25441_not ; n25594
g25339 and n25302_not n25594_not ; n25595
g25340 and n25593 n25595_not ; n25596
g25341 and n25593_not n25595 ; n25597
g25342 and n25596_not n25597_not ; n25598
g25343 and n25451_not n25598 ; n25599
g25344 and n25451 n25598_not ; n25600
g25345 and n25599_not n25600_not ; f[105]
g25346 and n25567_not n25573_not ; n25602
g25347 and b[62] n6902 ; n25603
g25348 and b[63] n6590 ; n25604
g25349 and n25603_not n25604_not ; n25605
g25350 and n6598_not n25605 ; n25606
g25351 and n13800 n25605 ; n25607
g25352 and n25606_not n25607_not ; n25608
g25353 and a[44] n25608_not ; n25609
g25354 and a[44]_not n25608 ; n25610
g25355 and n25609_not n25610_not ; n25611
g25356 and n25602_not n25611_not ; n25612
g25357 and n25602 n25611 ; n25613
g25358 and n25612_not n25613_not ; n25614
g25359 and b[61] n7446 ; n25615
g25360 and b[59] n7787 ; n25616
g25361 and b[60] n7441 ; n25617
g25362 and n25616_not n25617_not ; n25618
g25363 and n25615_not n25618 ; n25619
g25364 and n7449 n12969 ; n25620
g25365 and n25619 n25620_not ; n25621
g25366 and a[47] n25621_not ; n25622
g25367 and a[47] n25622_not ; n25623
g25368 and n25621_not n25622_not ; n25624
g25369 and n25623_not n25624_not ; n25625
g25370 and n25562_not n25564_not ; n25626
g25371 and n25556_not n25558_not ; n25627
g25372 and n25508_not n25514_not ; n25628
g25373 and b[42] n13903 ; n25629
g25374 and b[43] n13488_not ; n25630
g25375 and n25629_not n25630_not ; n25631
g25376 and a[41]_not n25146_not ; n25632
g25377 and n25495_not n25632_not ; n25633
g25378 and n25631 n25633_not ; n25634
g25379 and n25631 n25634_not ; n25635
g25380 and n25633_not n25634_not ; n25636
g25381 and n25635_not n25636_not ; n25637
g25382 and b[46] n12668 ; n25638
g25383 and b[44] n13047 ; n25639
g25384 and b[45] n12663 ; n25640
g25385 and n25639_not n25640_not ; n25641
g25386 and n25638_not n25641 ; n25642
g25387 and n12671_not n25642 ; n25643
g25388 and n7677_not n25642 ; n25644
g25389 and n25643_not n25644_not ; n25645
g25390 and a[62] n25645_not ; n25646
g25391 and a[62]_not n25645 ; n25647
g25392 and n25646_not n25647_not ; n25648
g25393 and n25637_not n25648_not ; n25649
g25394 and n25637 n25648 ; n25650
g25395 and n25649_not n25650_not ; n25651
g25396 and n25628_not n25651 ; n25652
g25397 and n25628 n25651_not ; n25653
g25398 and n25652_not n25653_not ; n25654
g25399 and b[49] n11531 ; n25655
g25400 and b[47] n11896 ; n25656
g25401 and b[48] n11526 ; n25657
g25402 and n25656_not n25657_not ; n25658
g25403 and n25655_not n25658 ; n25659
g25404 and n8625 n11534 ; n25660
g25405 and n25659 n25660_not ; n25661
g25406 and a[59] n25661_not ; n25662
g25407 and a[59] n25662_not ; n25663
g25408 and n25661_not n25662_not ; n25664
g25409 and n25663_not n25664_not ; n25665
g25410 and n25654 n25665_not ; n25666
g25411 and n25654 n25666_not ; n25667
g25412 and n25665_not n25666_not ; n25668
g25413 and n25667_not n25668_not ; n25669
g25414 and n25527_not n25533_not ; n25670
g25415 and n25669 n25670 ; n25671
g25416 and n25669_not n25670_not ; n25672
g25417 and n25671_not n25672_not ; n25673
g25418 and b[52] n10426 ; n25674
g25419 and b[50] n10796 ; n25675
g25420 and b[51] n10421 ; n25676
g25421 and n25675_not n25676_not ; n25677
g25422 and n25674_not n25677 ; n25678
g25423 and n9628 n10429 ; n25679
g25424 and n25678 n25679_not ; n25680
g25425 and a[56] n25680_not ; n25681
g25426 and a[56] n25681_not ; n25682
g25427 and n25680_not n25681_not ; n25683
g25428 and n25682_not n25683_not ; n25684
g25429 and n25673 n25684_not ; n25685
g25430 and n25673 n25685_not ; n25686
g25431 and n25684_not n25685_not ; n25687
g25432 and n25686_not n25687_not ; n25688
g25433 and n25536_not n25540_not ; n25689
g25434 and n25688 n25689 ; n25690
g25435 and n25688_not n25689_not ; n25691
g25436 and n25690_not n25691_not ; n25692
g25437 and b[55] n9339 ; n25693
g25438 and b[53] n9732 ; n25694
g25439 and b[54] n9334 ; n25695
g25440 and n25694_not n25695_not ; n25696
g25441 and n25693_not n25696 ; n25697
g25442 and n9342 n10684 ; n25698
g25443 and n25697 n25698_not ; n25699
g25444 and a[53] n25699_not ; n25700
g25445 and a[53] n25700_not ; n25701
g25446 and n25699_not n25700_not ; n25702
g25447 and n25701_not n25702_not ; n25703
g25448 and n25692 n25703_not ; n25704
g25449 and n25692 n25704_not ; n25705
g25450 and n25703_not n25704_not ; n25706
g25451 and n25705_not n25706_not ; n25707
g25452 and n25627_not n25707 ; n25708
g25453 and n25627 n25707_not ; n25709
g25454 and n25708_not n25709_not ; n25710
g25455 and b[58] n8362 ; n25711
g25456 and b[56] n8715 ; n25712
g25457 and b[57] n8357 ; n25713
g25458 and n25712_not n25713_not ; n25714
g25459 and n25711_not n25714 ; n25715
g25460 and n8365 n11436 ; n25716
g25461 and n25715 n25716_not ; n25717
g25462 and a[50] n25717_not ; n25718
g25463 and a[50] n25718_not ; n25719
g25464 and n25717_not n25718_not ; n25720
g25465 and n25719_not n25720_not ; n25721
g25466 and n25710 n25721 ; n25722
g25467 and n25710_not n25721_not ; n25723
g25468 and n25722_not n25723_not ; n25724
g25469 and n25626_not n25724 ; n25725
g25470 and n25626_not n25725_not ; n25726
g25471 and n25724 n25725_not ; n25727
g25472 and n25726_not n25727_not ; n25728
g25473 and n25625_not n25728_not ; n25729
g25474 and n25625_not n25729_not ; n25730
g25475 and n25728_not n25729_not ; n25731
g25476 and n25730_not n25731_not ; n25732
g25477 and n25614 n25732_not ; n25733
g25478 and n25614 n25733_not ; n25734
g25479 and n25732_not n25733_not ; n25735
g25480 and n25734_not n25735_not ; n25736
g25481 and n25586_not n25592_not ; n25737
g25482 and n25736 n25737 ; n25738
g25483 and n25736_not n25737_not ; n25739
g25484 and n25738_not n25739_not ; n25740
g25485 and n25596_not n25599_not ; n25741
g25486 and n25740 n25741_not ; n25742
g25487 and n25740_not n25741 ; n25743
g25488 and n25742_not n25743_not ; f[106]
g25489 and n25739_not n25742_not ; n25745
g25490 and n25612_not n25733_not ; n25746
g25491 and n25725_not n25729_not ; n25747
g25492 and b[63] n6902 ; n25748
g25493 and n6598 n13797 ; n25749
g25494 and n25748_not n25749_not ; n25750
g25495 and a[44] n25750_not ; n25751
g25496 and a[44] n25751_not ; n25752
g25497 and n25750_not n25751_not ; n25753
g25498 and n25752_not n25753_not ; n25754
g25499 and n25747_not n25754_not ; n25755
g25500 and n25747_not n25755_not ; n25756
g25501 and n25754_not n25755_not ; n25757
g25502 and n25756_not n25757_not ; n25758
g25503 and b[59] n8362 ; n25759
g25504 and b[57] n8715 ; n25760
g25505 and b[58] n8357 ; n25761
g25506 and n25760_not n25761_not ; n25762
g25507 and n25759_not n25762 ; n25763
g25508 and n8365 n12179 ; n25764
g25509 and n25763 n25764_not ; n25765
g25510 and a[50] n25765_not ; n25766
g25511 and a[50] n25766_not ; n25767
g25512 and n25765_not n25766_not ; n25768
g25513 and n25767_not n25768_not ; n25769
g25514 and n25691_not n25704_not ; n25770
g25515 and b[56] n9339 ; n25771
g25516 and b[54] n9732 ; n25772
g25517 and b[55] n9334 ; n25773
g25518 and n25772_not n25773_not ; n25774
g25519 and n25771_not n25774 ; n25775
g25520 and n9342 n10708 ; n25776
g25521 and n25775 n25776_not ; n25777
g25522 and a[53] n25777_not ; n25778
g25523 and a[53] n25778_not ; n25779
g25524 and n25777_not n25778_not ; n25780
g25525 and n25779_not n25780_not ; n25781
g25526 and n25672_not n25685_not ; n25782
g25527 and b[53] n10426 ; n25783
g25528 and b[51] n10796 ; n25784
g25529 and b[52] n10421 ; n25785
g25530 and n25784_not n25785_not ; n25786
g25531 and n25783_not n25786 ; n25787
g25532 and n9972 n10429 ; n25788
g25533 and n25787 n25788_not ; n25789
g25534 and a[56] n25789_not ; n25790
g25535 and a[56] n25790_not ; n25791
g25536 and n25789_not n25790_not ; n25792
g25537 and n25791_not n25792_not ; n25793
g25538 and n25652_not n25666_not ; n25794
g25539 and b[50] n11531 ; n25795
g25540 and b[48] n11896 ; n25796
g25541 and b[49] n11526 ; n25797
g25542 and n25796_not n25797_not ; n25798
g25543 and n25795_not n25798 ; n25799
g25544 and n8949 n11534 ; n25800
g25545 and n25799 n25800_not ; n25801
g25546 and a[59] n25801_not ; n25802
g25547 and a[59] n25802_not ; n25803
g25548 and n25801_not n25802_not ; n25804
g25549 and n25803_not n25804_not ; n25805
g25550 and n25634_not n25649_not ; n25806
g25551 and b[43] n13903 ; n25807
g25552 and b[44] n13488_not ; n25808
g25553 and n25807_not n25808_not ; n25809
g25554 and n25631 n25809_not ; n25810
g25555 and n25631_not n25809 ; n25811
g25556 and n25810_not n25811_not ; n25812
g25557 and b[47] n12668 ; n25813
g25558 and b[45] n13047 ; n25814
g25559 and b[46] n12663 ; n25815
g25560 and n25814_not n25815_not ; n25816
g25561 and n25813_not n25816 ; n25817
g25562 and n12671_not n25817 ; n25818
g25563 and n7703_not n25817 ; n25819
g25564 and n25818_not n25819_not ; n25820
g25565 and a[62] n25820_not ; n25821
g25566 and a[62]_not n25820 ; n25822
g25567 and n25821_not n25822_not ; n25823
g25568 and n25812 n25823_not ; n25824
g25569 and n25812_not n25823 ; n25825
g25570 and n25824_not n25825_not ; n25826
g25571 and n25806_not n25826 ; n25827
g25572 and n25806_not n25827_not ; n25828
g25573 and n25826 n25827_not ; n25829
g25574 and n25828_not n25829_not ; n25830
g25575 and n25805_not n25830_not ; n25831
g25576 and n25805 n25829_not ; n25832
g25577 and n25828_not n25832 ; n25833
g25578 and n25831_not n25833_not ; n25834
g25579 and n25794_not n25834 ; n25835
g25580 and n25794_not n25835_not ; n25836
g25581 and n25834 n25835_not ; n25837
g25582 and n25836_not n25837_not ; n25838
g25583 and n25793_not n25838_not ; n25839
g25584 and n25793 n25837_not ; n25840
g25585 and n25836_not n25840 ; n25841
g25586 and n25839_not n25841_not ; n25842
g25587 and n25782_not n25842 ; n25843
g25588 and n25782_not n25843_not ; n25844
g25589 and n25842 n25843_not ; n25845
g25590 and n25844_not n25845_not ; n25846
g25591 and n25781_not n25846_not ; n25847
g25592 and n25781 n25845_not ; n25848
g25593 and n25844_not n25848 ; n25849
g25594 and n25847_not n25849_not ; n25850
g25595 and n25770_not n25850 ; n25851
g25596 and n25770 n25850_not ; n25852
g25597 and n25851_not n25852_not ; n25853
g25598 and n25769_not n25853 ; n25854
g25599 and n25853 n25854_not ; n25855
g25600 and n25769_not n25854_not ; n25856
g25601 and n25855_not n25856_not ; n25857
g25602 and n25627_not n25707_not ; n25858
g25603 and n25723_not n25858_not ; n25859
g25604 and n25857_not n25859_not ; n25860
g25605 and n25857_not n25860_not ; n25861
g25606 and n25859_not n25860_not ; n25862
g25607 and n25861_not n25862_not ; n25863
g25608 and b[62] n7446 ; n25864
g25609 and b[60] n7787 ; n25865
g25610 and b[61] n7441 ; n25866
g25611 and n25865_not n25866_not ; n25867
g25612 and n25864_not n25867 ; n25868
g25613 and n7449 n13370 ; n25869
g25614 and n25868 n25869_not ; n25870
g25615 and a[47] n25870_not ; n25871
g25616 and a[47] n25871_not ; n25872
g25617 and n25870_not n25871_not ; n25873
g25618 and n25872_not n25873_not ; n25874
g25619 and n25863_not n25874_not ; n25875
g25620 and n25863_not n25875_not ; n25876
g25621 and n25874_not n25875_not ; n25877
g25622 and n25876_not n25877_not ; n25878
g25623 and n25758_not n25878 ; n25879
g25624 and n25758 n25878_not ; n25880
g25625 and n25879_not n25880_not ; n25881
g25626 and n25746_not n25881_not ; n25882
g25627 and n25746 n25881 ; n25883
g25628 and n25882_not n25883_not ; n25884
g25629 and n25745_not n25884 ; n25885
g25630 and n25745 n25884_not ; n25886
g25631 and n25885_not n25886_not ; f[107]
g25632 and n25882_not n25885_not ; n25888
g25633 and b[63] n7446 ; n25889
g25634 and b[61] n7787 ; n25890
g25635 and b[62] n7441 ; n25891
g25636 and n25890_not n25891_not ; n25892
g25637 and n25889_not n25892 ; n25893
g25638 and n7449 n13771 ; n25894
g25639 and n25893 n25894_not ; n25895
g25640 and a[47] n25895_not ; n25896
g25641 and a[47] n25896_not ; n25897
g25642 and n25895_not n25896_not ; n25898
g25643 and n25897_not n25898_not ; n25899
g25644 and n25851_not n25854_not ; n25900
g25645 and b[60] n8362 ; n25901
g25646 and b[58] n8715 ; n25902
g25647 and b[59] n8357 ; n25903
g25648 and n25902_not n25903_not ; n25904
g25649 and n25901_not n25904 ; n25905
g25650 and n8365 n12211 ; n25906
g25651 and n25905 n25906_not ; n25907
g25652 and a[50] n25907_not ; n25908
g25653 and a[50] n25908_not ; n25909
g25654 and n25907_not n25908_not ; n25910
g25655 and n25909_not n25910_not ; n25911
g25656 and n25843_not n25847_not ; n25912
g25657 and b[57] n9339 ; n25913
g25658 and b[55] n9732 ; n25914
g25659 and b[56] n9334 ; n25915
g25660 and n25914_not n25915_not ; n25916
g25661 and n25913_not n25916 ; n25917
g25662 and n9342 n11410 ; n25918
g25663 and n25917 n25918_not ; n25919
g25664 and a[53] n25919_not ; n25920
g25665 and a[53] n25920_not ; n25921
g25666 and n25919_not n25920_not ; n25922
g25667 and n25921_not n25922_not ; n25923
g25668 and n25835_not n25839_not ; n25924
g25669 and b[54] n10426 ; n25925
g25670 and b[52] n10796 ; n25926
g25671 and b[53] n10421 ; n25927
g25672 and n25926_not n25927_not ; n25928
g25673 and n25925_not n25928 ; n25929
g25674 and n9998 n10429 ; n25930
g25675 and n25929 n25930_not ; n25931
g25676 and a[56] n25931_not ; n25932
g25677 and a[56] n25932_not ; n25933
g25678 and n25931_not n25932_not ; n25934
g25679 and n25933_not n25934_not ; n25935
g25680 and n25827_not n25831_not ; n25936
g25681 and n25810_not n25824_not ; n25937
g25682 and b[44] n13903 ; n25938
g25683 and b[45] n13488_not ; n25939
g25684 and n25938_not n25939_not ; n25940
g25685 and a[44]_not n25940_not ; n25941
g25686 and a[44] n25940 ; n25942
g25687 and n25941_not n25942_not ; n25943
g25688 and n25631_not n25943 ; n25944
g25689 and n25631_not n25944_not ; n25945
g25690 and n25943 n25944_not ; n25946
g25691 and n25945_not n25946_not ; n25947
g25692 and n25937_not n25947_not ; n25948
g25693 and n25937_not n25948_not ; n25949
g25694 and n25947_not n25948_not ; n25950
g25695 and n25949_not n25950_not ; n25951
g25696 and b[48] n12668 ; n25952
g25697 and b[46] n13047 ; n25953
g25698 and b[47] n12663 ; n25954
g25699 and n25953_not n25954_not ; n25955
g25700 and n25952_not n25955 ; n25956
g25701 and n8009 n12671 ; n25957
g25702 and n25956 n25957_not ; n25958
g25703 and a[62] n25958_not ; n25959
g25704 and a[62] n25959_not ; n25960
g25705 and n25958_not n25959_not ; n25961
g25706 and n25960_not n25961_not ; n25962
g25707 and n25951_not n25962_not ; n25963
g25708 and n25951_not n25963_not ; n25964
g25709 and n25962_not n25963_not ; n25965
g25710 and n25964_not n25965_not ; n25966
g25711 and b[51] n11531 ; n25967
g25712 and b[49] n11896 ; n25968
g25713 and b[50] n11526 ; n25969
g25714 and n25968_not n25969_not ; n25970
g25715 and n25967_not n25970 ; n25971
g25716 and n8976 n11534 ; n25972
g25717 and n25971 n25972_not ; n25973
g25718 and a[59] n25973_not ; n25974
g25719 and a[59] n25974_not ; n25975
g25720 and n25973_not n25974_not ; n25976
g25721 and n25975_not n25976_not ; n25977
g25722 and n25966 n25977 ; n25978
g25723 and n25966_not n25977_not ; n25979
g25724 and n25978_not n25979_not ; n25980
g25725 and n25936_not n25980 ; n25981
g25726 and n25936 n25980_not ; n25982
g25727 and n25981_not n25982_not ; n25983
g25728 and n25935 n25983_not ; n25984
g25729 and n25935_not n25983 ; n25985
g25730 and n25984_not n25985_not ; n25986
g25731 and n25924_not n25986 ; n25987
g25732 and n25924 n25986_not ; n25988
g25733 and n25987_not n25988_not ; n25989
g25734 and n25923 n25989_not ; n25990
g25735 and n25923_not n25989 ; n25991
g25736 and n25990_not n25991_not ; n25992
g25737 and n25912_not n25992 ; n25993
g25738 and n25912 n25992_not ; n25994
g25739 and n25993_not n25994_not ; n25995
g25740 and n25911 n25995_not ; n25996
g25741 and n25911_not n25995 ; n25997
g25742 and n25996_not n25997_not ; n25998
g25743 and n25900_not n25998 ; n25999
g25744 and n25900 n25998_not ; n26000
g25745 and n25999_not n26000_not ; n26001
g25746 and n25899_not n26001 ; n26002
g25747 and n26001 n26002_not ; n26003
g25748 and n25899_not n26002_not ; n26004
g25749 and n26003_not n26004_not ; n26005
g25750 and n25860_not n25875_not ; n26006
g25751 and n26005 n26006 ; n26007
g25752 and n26005_not n26006_not ; n26008
g25753 and n26007_not n26008_not ; n26009
g25754 and n25758_not n25878_not ; n26010
g25755 and n25755_not n26010_not ; n26011
g25756 and n26009 n26011_not ; n26012
g25757 and n26009_not n26011 ; n26013
g25758 and n26012_not n26013_not ; n26014
g25759 and n25888_not n26014 ; n26015
g25760 and n25888 n26014_not ; n26016
g25761 and n26015_not n26016_not ; f[108]
g25762 and n25997_not n25999_not ; n26018
g25763 and b[62] n7787 ; n26019
g25764 and b[63] n7441 ; n26020
g25765 and n26019_not n26020_not ; n26021
g25766 and n7449_not n26021 ; n26022
g25767 and n13800 n26021 ; n26023
g25768 and n26022_not n26023_not ; n26024
g25769 and a[47] n26024_not ; n26025
g25770 and a[47]_not n26024 ; n26026
g25771 and n26025_not n26026_not ; n26027
g25772 and n26018_not n26027_not ; n26028
g25773 and n26018 n26027 ; n26029
g25774 and n26028_not n26029_not ; n26030
g25775 and b[61] n8362 ; n26031
g25776 and b[59] n8715 ; n26032
g25777 and b[60] n8357 ; n26033
g25778 and n26032_not n26033_not ; n26034
g25779 and n26031_not n26034 ; n26035
g25780 and n8365 n12969 ; n26036
g25781 and n26035 n26036_not ; n26037
g25782 and a[50] n26037_not ; n26038
g25783 and a[50] n26038_not ; n26039
g25784 and n26037_not n26038_not ; n26040
g25785 and n26039_not n26040_not ; n26041
g25786 and n25991_not n25993_not ; n26042
g25787 and n25985_not n25987_not ; n26043
g25788 and b[55] n10426 ; n26044
g25789 and b[53] n10796 ; n26045
g25790 and b[54] n10421 ; n26046
g25791 and n26045_not n26046_not ; n26047
g25792 and n26044_not n26047 ; n26048
g25793 and n10429 n10684 ; n26049
g25794 and n26048 n26049_not ; n26050
g25795 and a[56] n26050_not ; n26051
g25796 and a[56] n26051_not ; n26052
g25797 and n26050_not n26051_not ; n26053
g25798 and n26052_not n26053_not ; n26054
g25799 and n25979_not n25981_not ; n26055
g25800 and b[52] n11531 ; n26056
g25801 and b[50] n11896 ; n26057
g25802 and b[51] n11526 ; n26058
g25803 and n26057_not n26058_not ; n26059
g25804 and n26056_not n26059 ; n26060
g25805 and n9628 n11534 ; n26061
g25806 and n26060 n26061_not ; n26062
g25807 and a[59] n26062_not ; n26063
g25808 and a[59] n26063_not ; n26064
g25809 and n26062_not n26063_not ; n26065
g25810 and n26064_not n26065_not ; n26066
g25811 and n25948_not n25963_not ; n26067
g25812 and b[45] n13903 ; n26068
g25813 and b[46] n13488_not ; n26069
g25814 and n26068_not n26069_not ; n26070
g25815 and n25941_not n25944_not ; n26071
g25816 and n26070_not n26071 ; n26072
g25817 and n26070 n26071_not ; n26073
g25818 and n26072_not n26073_not ; n26074
g25819 and b[49] n12668 ; n26075
g25820 and b[47] n13047 ; n26076
g25821 and b[48] n12663 ; n26077
g25822 and n26076_not n26077_not ; n26078
g25823 and n26075_not n26078 ; n26079
g25824 and n8625 n12671 ; n26080
g25825 and n26079 n26080_not ; n26081
g25826 and a[62] n26081_not ; n26082
g25827 and a[62] n26082_not ; n26083
g25828 and n26081_not n26082_not ; n26084
g25829 and n26083_not n26084_not ; n26085
g25830 and n26074_not n26085 ; n26086
g25831 and n26074 n26085_not ; n26087
g25832 and n26086_not n26087_not ; n26088
g25833 and n26067_not n26088 ; n26089
g25834 and n26067_not n26089_not ; n26090
g25835 and n26088 n26089_not ; n26091
g25836 and n26090_not n26091_not ; n26092
g25837 and n26066_not n26092_not ; n26093
g25838 and n26066 n26091_not ; n26094
g25839 and n26090_not n26094 ; n26095
g25840 and n26093_not n26095_not ; n26096
g25841 and n26055_not n26096 ; n26097
g25842 and n26055 n26096_not ; n26098
g25843 and n26097_not n26098_not ; n26099
g25844 and n26054_not n26099 ; n26100
g25845 and n26099 n26100_not ; n26101
g25846 and n26054_not n26100_not ; n26102
g25847 and n26101_not n26102_not ; n26103
g25848 and n26043_not n26103 ; n26104
g25849 and n26043 n26103_not ; n26105
g25850 and n26104_not n26105_not ; n26106
g25851 and b[58] n9339 ; n26107
g25852 and b[56] n9732 ; n26108
g25853 and b[57] n9334 ; n26109
g25854 and n26108_not n26109_not ; n26110
g25855 and n26107_not n26110 ; n26111
g25856 and n9342 n11436 ; n26112
g25857 and n26111 n26112_not ; n26113
g25858 and a[53] n26113_not ; n26114
g25859 and a[53] n26114_not ; n26115
g25860 and n26113_not n26114_not ; n26116
g25861 and n26115_not n26116_not ; n26117
g25862 and n26106 n26117 ; n26118
g25863 and n26106_not n26117_not ; n26119
g25864 and n26118_not n26119_not ; n26120
g25865 and n26042_not n26120 ; n26121
g25866 and n26042_not n26121_not ; n26122
g25867 and n26120 n26121_not ; n26123
g25868 and n26122_not n26123_not ; n26124
g25869 and n26041_not n26124_not ; n26125
g25870 and n26041_not n26125_not ; n26126
g25871 and n26124_not n26125_not ; n26127
g25872 and n26126_not n26127_not ; n26128
g25873 and n26030 n26128_not ; n26129
g25874 and n26030 n26129_not ; n26130
g25875 and n26128_not n26129_not ; n26131
g25876 and n26130_not n26131_not ; n26132
g25877 and n26002_not n26008_not ; n26133
g25878 and n26132 n26133 ; n26134
g25879 and n26132_not n26133_not ; n26135
g25880 and n26134_not n26135_not ; n26136
g25881 and n26012_not n26015_not ; n26137
g25882 and n26136 n26137_not ; n26138
g25883 and n26136_not n26137 ; n26139
g25884 and n26138_not n26139_not ; f[109]
g25885 and b[59] n9339 ; n26141
g25886 and b[57] n9732 ; n26142
g25887 and b[58] n9334 ; n26143
g25888 and n26142_not n26143_not ; n26144
g25889 and n26141_not n26144 ; n26145
g25890 and n9342 n12179 ; n26146
g25891 and n26145 n26146_not ; n26147
g25892 and a[53] n26147_not ; n26148
g25893 and a[53] n26148_not ; n26149
g25894 and n26147_not n26148_not ; n26150
g25895 and n26149_not n26150_not ; n26151
g25896 and n26097_not n26100_not ; n26152
g25897 and b[56] n10426 ; n26153
g25898 and b[54] n10796 ; n26154
g25899 and b[55] n10421 ; n26155
g25900 and n26154_not n26155_not ; n26156
g25901 and n26153_not n26156 ; n26157
g25902 and n10429 n10708 ; n26158
g25903 and n26157 n26158_not ; n26159
g25904 and a[56] n26159_not ; n26160
g25905 and a[56] n26160_not ; n26161
g25906 and n26159_not n26160_not ; n26162
g25907 and n26161_not n26162_not ; n26163
g25908 and n26089_not n26093_not ; n26164
g25909 and b[53] n11531 ; n26165
g25910 and b[51] n11896 ; n26166
g25911 and b[52] n11526 ; n26167
g25912 and n26166_not n26167_not ; n26168
g25913 and n26165_not n26168 ; n26169
g25914 and n9972 n11534 ; n26170
g25915 and n26169 n26170_not ; n26171
g25916 and a[59] n26171_not ; n26172
g25917 and a[59] n26172_not ; n26173
g25918 and n26171_not n26172_not ; n26174
g25919 and n26173_not n26174_not ; n26175
g25920 and n26073_not n26087_not ; n26176
g25921 and b[46] n13903 ; n26177
g25922 and b[47] n13488_not ; n26178
g25923 and n26177_not n26178_not ; n26179
g25924 and n26070 n26179_not ; n26180
g25925 and n26070_not n26179 ; n26181
g25926 and n26176_not n26181_not ; n26182
g25927 and n26180_not n26182 ; n26183
g25928 and n26176_not n26183_not ; n26184
g25929 and n26181_not n26183_not ; n26185
g25930 and n26180_not n26185 ; n26186
g25931 and n26184_not n26186_not ; n26187
g25932 and b[50] n12668 ; n26188
g25933 and b[48] n13047 ; n26189
g25934 and b[49] n12663 ; n26190
g25935 and n26189_not n26190_not ; n26191
g25936 and n26188_not n26191 ; n26192
g25937 and n8949 n12671 ; n26193
g25938 and n26192 n26193_not ; n26194
g25939 and a[62] n26194_not ; n26195
g25940 and a[62] n26195_not ; n26196
g25941 and n26194_not n26195_not ; n26197
g25942 and n26196_not n26197_not ; n26198
g25943 and n26187_not n26198 ; n26199
g25944 and n26187 n26198_not ; n26200
g25945 and n26199_not n26200_not ; n26201
g25946 and n26175_not n26201_not ; n26202
g25947 and n26175 n26201 ; n26203
g25948 and n26202_not n26203_not ; n26204
g25949 and n26164_not n26204 ; n26205
g25950 and n26164_not n26205_not ; n26206
g25951 and n26204 n26205_not ; n26207
g25952 and n26206_not n26207_not ; n26208
g25953 and n26163_not n26208_not ; n26209
g25954 and n26163 n26207_not ; n26210
g25955 and n26206_not n26210 ; n26211
g25956 and n26209_not n26211_not ; n26212
g25957 and n26152_not n26212 ; n26213
g25958 and n26152 n26212_not ; n26214
g25959 and n26213_not n26214_not ; n26215
g25960 and n26151_not n26215 ; n26216
g25961 and n26215 n26216_not ; n26217
g25962 and n26151_not n26216_not ; n26218
g25963 and n26217_not n26218_not ; n26219
g25964 and n26043_not n26103_not ; n26220
g25965 and n26119_not n26220_not ; n26221
g25966 and n26219_not n26221_not ; n26222
g25967 and n26219_not n26222_not ; n26223
g25968 and n26221_not n26222_not ; n26224
g25969 and n26223_not n26224_not ; n26225
g25970 and b[62] n8362 ; n26226
g25971 and b[60] n8715 ; n26227
g25972 and b[61] n8357 ; n26228
g25973 and n26227_not n26228_not ; n26229
g25974 and n26226_not n26229 ; n26230
g25975 and n8365 n13370 ; n26231
g25976 and n26230 n26231_not ; n26232
g25977 and a[50] n26232_not ; n26233
g25978 and a[50] n26233_not ; n26234
g25979 and n26232_not n26233_not ; n26235
g25980 and n26234_not n26235_not ; n26236
g25981 and n26225_not n26236_not ; n26237
g25982 and n26225_not n26237_not ; n26238
g25983 and n26236_not n26237_not ; n26239
g25984 and n26238_not n26239_not ; n26240
g25985 and n26121_not n26125_not ; n26241
g25986 and b[63] n7787 ; n26242
g25987 and n7449_not n26242_not ; n26243
g25988 and n13797_not n26242_not ; n26244
g25989 and n26243_not n26244_not ; n26245
g25990 and a[47] n26245_not ; n26246
g25991 and a[47]_not n26245 ; n26247
g25992 and n26246_not n26247_not ; n26248
g25993 and n26241_not n26248_not ; n26249
g25994 and n26241 n26248 ; n26250
g25995 and n26249_not n26250_not ; n26251
g25996 and n26240_not n26251 ; n26252
g25997 and n26240_not n26252_not ; n26253
g25998 and n26251 n26252_not ; n26254
g25999 and n26253_not n26254_not ; n26255
g26000 and n26028_not n26129_not ; n26256
g26001 and n26255 n26256 ; n26257
g26002 and n26255_not n26256_not ; n26258
g26003 and n26257_not n26258_not ; n26259
g26004 and n26135_not n26138_not ; n26260
g26005 and n26259 n26260_not ; n26261
g26006 and n26259_not n26260 ; n26262
g26007 and n26261_not n26262_not ; f[110]
g26008 and b[63] n8362 ; n26264
g26009 and b[61] n8715 ; n26265
g26010 and b[62] n8357 ; n26266
g26011 and n26265_not n26266_not ; n26267
g26012 and n26264_not n26267 ; n26268
g26013 and n8365 n13771 ; n26269
g26014 and n26268 n26269_not ; n26270
g26015 and a[50] n26270_not ; n26271
g26016 and a[50] n26271_not ; n26272
g26017 and n26270_not n26271_not ; n26273
g26018 and n26272_not n26273_not ; n26274
g26019 and n26213_not n26216_not ; n26275
g26020 and b[60] n9339 ; n26276
g26021 and b[58] n9732 ; n26277
g26022 and b[59] n9334 ; n26278
g26023 and n26277_not n26278_not ; n26279
g26024 and n26276_not n26279 ; n26280
g26025 and n9342 n12211 ; n26281
g26026 and n26280 n26281_not ; n26282
g26027 and a[53] n26282_not ; n26283
g26028 and a[53] n26283_not ; n26284
g26029 and n26282_not n26283_not ; n26285
g26030 and n26284_not n26285_not ; n26286
g26031 and n26205_not n26209_not ; n26287
g26032 and b[57] n10426 ; n26288
g26033 and b[55] n10796 ; n26289
g26034 and b[56] n10421 ; n26290
g26035 and n26289_not n26290_not ; n26291
g26036 and n26288_not n26291 ; n26292
g26037 and n10429 n11410 ; n26293
g26038 and n26292 n26293_not ; n26294
g26039 and a[56] n26294_not ; n26295
g26040 and a[56] n26295_not ; n26296
g26041 and n26294_not n26295_not ; n26297
g26042 and n26296_not n26297_not ; n26298
g26043 and n26187_not n26198_not ; n26299
g26044 and n26202_not n26299_not ; n26300
g26045 and b[51] n12668 ; n26301
g26046 and b[49] n13047 ; n26302
g26047 and b[50] n12663 ; n26303
g26048 and n26302_not n26303_not ; n26304
g26049 and n26301_not n26304 ; n26305
g26050 and n8976 n12671 ; n26306
g26051 and n26305 n26306_not ; n26307
g26052 and a[62] n26307_not ; n26308
g26053 and a[62] n26308_not ; n26309
g26054 and n26307_not n26308_not ; n26310
g26055 and n26309_not n26310_not ; n26311
g26056 and b[47] n13903 ; n26312
g26057 and b[48] n13488_not ; n26313
g26058 and n26312_not n26313_not ; n26314
g26059 and a[47] n26179_not ; n26315
g26060 and a[47]_not n26179 ; n26316
g26061 and n26315_not n26316_not ; n26317
g26062 and n26314_not n26317_not ; n26318
g26063 and n26314 n26317 ; n26319
g26064 and n26318_not n26319_not ; n26320
g26065 and n26311_not n26320 ; n26321
g26066 and n26311_not n26321_not ; n26322
g26067 and n26320 n26321_not ; n26323
g26068 and n26322_not n26323_not ; n26324
g26069 and n26185_not n26324_not ; n26325
g26070 and n26185_not n26325_not ; n26326
g26071 and n26324_not n26325_not ; n26327
g26072 and n26326_not n26327_not ; n26328
g26073 and b[54] n11531 ; n26329
g26074 and b[52] n11896 ; n26330
g26075 and b[53] n11526 ; n26331
g26076 and n26330_not n26331_not ; n26332
g26077 and n26329_not n26332 ; n26333
g26078 and n9998 n11534 ; n26334
g26079 and n26333 n26334_not ; n26335
g26080 and a[59] n26335_not ; n26336
g26081 and a[59] n26336_not ; n26337
g26082 and n26335_not n26336_not ; n26338
g26083 and n26337_not n26338_not ; n26339
g26084 and n26328 n26339 ; n26340
g26085 and n26328_not n26339_not ; n26341
g26086 and n26340_not n26341_not ; n26342
g26087 and n26300_not n26342 ; n26343
g26088 and n26300 n26342_not ; n26344
g26089 and n26343_not n26344_not ; n26345
g26090 and n26298 n26345_not ; n26346
g26091 and n26298_not n26345 ; n26347
g26092 and n26346_not n26347_not ; n26348
g26093 and n26287_not n26348 ; n26349
g26094 and n26287 n26348_not ; n26350
g26095 and n26349_not n26350_not ; n26351
g26096 and n26286 n26351_not ; n26352
g26097 and n26286_not n26351 ; n26353
g26098 and n26352_not n26353_not ; n26354
g26099 and n26275_not n26354 ; n26355
g26100 and n26275 n26354_not ; n26356
g26101 and n26355_not n26356_not ; n26357
g26102 and n26274_not n26357 ; n26358
g26103 and n26357 n26358_not ; n26359
g26104 and n26274_not n26358_not ; n26360
g26105 and n26359_not n26360_not ; n26361
g26106 and n26222_not n26237_not ; n26362
g26107 and n26361 n26362 ; n26363
g26108 and n26361_not n26362_not ; n26364
g26109 and n26363_not n26364_not ; n26365
g26110 and n26249_not n26252_not ; n26366
g26111 and n26365_not n26366 ; n26367
g26112 and n26365 n26366_not ; n26368
g26113 and n26367_not n26368_not ; n26369
g26114 and n26258_not n26261_not ; n26370
g26115 and n26369 n26370_not ; n26371
g26116 and n26369_not n26370 ; n26372
g26117 and n26371_not n26372_not ; f[111]
g26118 and b[62] n8715 ; n26374
g26119 and b[63] n8357 ; n26375
g26120 and n26374_not n26375_not ; n26376
g26121 and n8365 n13800_not ; n26377
g26122 and n26376 n26377_not ; n26378
g26123 and a[50] n26378_not ; n26379
g26124 and a[50] n26379_not ; n26380
g26125 and n26378_not n26379_not ; n26381
g26126 and n26380_not n26381_not ; n26382
g26127 and n26353_not n26355_not ; n26383
g26128 and b[61] n9339 ; n26384
g26129 and b[59] n9732 ; n26385
g26130 and b[60] n9334 ; n26386
g26131 and n26385_not n26386_not ; n26387
g26132 and n26384_not n26387 ; n26388
g26133 and n9342 n12969 ; n26389
g26134 and n26388 n26389_not ; n26390
g26135 and a[53] n26390_not ; n26391
g26136 and a[53] n26391_not ; n26392
g26137 and n26390_not n26391_not ; n26393
g26138 and n26392_not n26393_not ; n26394
g26139 and n26347_not n26349_not ; n26395
g26140 and b[58] n10426 ; n26396
g26141 and b[56] n10796 ; n26397
g26142 and b[57] n10421 ; n26398
g26143 and n26397_not n26398_not ; n26399
g26144 and n26396_not n26399 ; n26400
g26145 and n10429 n11436 ; n26401
g26146 and n26400 n26401_not ; n26402
g26147 and a[56] n26402_not ; n26403
g26148 and a[56] n26403_not ; n26404
g26149 and n26402_not n26403_not ; n26405
g26150 and n26404_not n26405_not ; n26406
g26151 and n26341_not n26343_not ; n26407
g26152 and b[55] n11531 ; n26408
g26153 and b[53] n11896 ; n26409
g26154 and b[54] n11526 ; n26410
g26155 and n26409_not n26410_not ; n26411
g26156 and n26408_not n26411 ; n26412
g26157 and n10684 n11534 ; n26413
g26158 and n26412 n26413_not ; n26414
g26159 and a[59] n26414_not ; n26415
g26160 and a[59] n26415_not ; n26416
g26161 and n26414_not n26415_not ; n26417
g26162 and n26416_not n26417_not ; n26418
g26163 and n26321_not n26325_not ; n26419
g26164 and b[48] n13903 ; n26420
g26165 and b[49] n13488_not ; n26421
g26166 and n26420_not n26421_not ; n26422
g26167 and a[47]_not n26179_not ; n26423
g26168 and n26318_not n26423_not ; n26424
g26169 and n26422 n26424_not ; n26425
g26170 and n26422_not n26424 ; n26426
g26171 and n26425_not n26426_not ; n26427
g26172 and b[52] n12668 ; n26428
g26173 and b[50] n13047 ; n26429
g26174 and b[51] n12663 ; n26430
g26175 and n26429_not n26430_not ; n26431
g26176 and n26428_not n26431 ; n26432
g26177 and n12671_not n26432 ; n26433
g26178 and n9628_not n26432 ; n26434
g26179 and n26433_not n26434_not ; n26435
g26180 and a[62] n26435_not ; n26436
g26181 and a[62]_not n26435 ; n26437
g26182 and n26436_not n26437_not ; n26438
g26183 and n26427 n26438_not ; n26439
g26184 and n26427_not n26438 ; n26440
g26185 and n26439_not n26440_not ; n26441
g26186 and n26419_not n26441 ; n26442
g26187 and n26419_not n26442_not ; n26443
g26188 and n26441 n26442_not ; n26444
g26189 and n26443_not n26444_not ; n26445
g26190 and n26418_not n26445_not ; n26446
g26191 and n26418 n26444_not ; n26447
g26192 and n26443_not n26447 ; n26448
g26193 and n26446_not n26448_not ; n26449
g26194 and n26407_not n26449 ; n26450
g26195 and n26407 n26449_not ; n26451
g26196 and n26450_not n26451_not ; n26452
g26197 and n26406_not n26452 ; n26453
g26198 and n26406 n26452_not ; n26454
g26199 and n26453_not n26454_not ; n26455
g26200 and n26395_not n26455 ; n26456
g26201 and n26395_not n26456_not ; n26457
g26202 and n26455 n26456_not ; n26458
g26203 and n26457_not n26458_not ; n26459
g26204 and n26394_not n26459_not ; n26460
g26205 and n26394 n26458_not ; n26461
g26206 and n26457_not n26461 ; n26462
g26207 and n26460_not n26462_not ; n26463
g26208 and n26383_not n26463 ; n26464
g26209 and n26383 n26463_not ; n26465
g26210 and n26464_not n26465_not ; n26466
g26211 and n26382_not n26466 ; n26467
g26212 and n26466 n26467_not ; n26468
g26213 and n26382_not n26467_not ; n26469
g26214 and n26468_not n26469_not ; n26470
g26215 and n26358_not n26364_not ; n26471
g26216 and n26470 n26471 ; n26472
g26217 and n26470_not n26471_not ; n26473
g26218 and n26472_not n26473_not ; n26474
g26219 and n26368_not n26371_not ; n26475
g26220 and n26474 n26475_not ; n26476
g26221 and n26474_not n26475 ; n26477
g26222 and n26476_not n26477_not ; f[112]
g26223 and b[59] n10426 ; n26479
g26224 and b[57] n10796 ; n26480
g26225 and b[58] n10421 ; n26481
g26226 and n26480_not n26481_not ; n26482
g26227 and n26479_not n26482 ; n26483
g26228 and n10429 n12179 ; n26484
g26229 and n26483 n26484_not ; n26485
g26230 and a[56] n26485_not ; n26486
g26231 and a[56] n26486_not ; n26487
g26232 and n26485_not n26486_not ; n26488
g26233 and n26487_not n26488_not ; n26489
g26234 and n26442_not n26446_not ; n26490
g26235 and b[53] n12668 ; n26491
g26236 and b[51] n13047 ; n26492
g26237 and b[52] n12663 ; n26493
g26238 and n26492_not n26493_not ; n26494
g26239 and n26491_not n26494 ; n26495
g26240 and n9972 n12671 ; n26496
g26241 and n26495 n26496_not ; n26497
g26242 and a[62] n26497_not ; n26498
g26243 and a[62] n26498_not ; n26499
g26244 and n26497_not n26498_not ; n26500
g26245 and n26499_not n26500_not ; n26501
g26246 and b[49] n13903 ; n26502
g26247 and b[50] n13488_not ; n26503
g26248 and n26502_not n26503_not ; n26504
g26249 and n26422 n26504_not ; n26505
g26250 and n26422 n26505_not ; n26506
g26251 and n26504_not n26505_not ; n26507
g26252 and n26506_not n26507_not ; n26508
g26253 and n26501_not n26508_not ; n26509
g26254 and n26501_not n26509_not ; n26510
g26255 and n26508_not n26509_not ; n26511
g26256 and n26510_not n26511_not ; n26512
g26257 and n26425_not n26439_not ; n26513
g26258 and n26512 n26513 ; n26514
g26259 and n26512_not n26513_not ; n26515
g26260 and n26514_not n26515_not ; n26516
g26261 and b[56] n11531 ; n26517
g26262 and b[54] n11896 ; n26518
g26263 and b[55] n11526 ; n26519
g26264 and n26518_not n26519_not ; n26520
g26265 and n26517_not n26520 ; n26521
g26266 and n10708 n11534 ; n26522
g26267 and n26521 n26522_not ; n26523
g26268 and a[59] n26523_not ; n26524
g26269 and a[59] n26524_not ; n26525
g26270 and n26523_not n26524_not ; n26526
g26271 and n26525_not n26526_not ; n26527
g26272 and n26516_not n26527 ; n26528
g26273 and n26516 n26527_not ; n26529
g26274 and n26528_not n26529_not ; n26530
g26275 and n26490_not n26530 ; n26531
g26276 and n26490 n26530_not ; n26532
g26277 and n26531_not n26532_not ; n26533
g26278 and n26489_not n26533 ; n26534
g26279 and n26533 n26534_not ; n26535
g26280 and n26489_not n26534_not ; n26536
g26281 and n26535_not n26536_not ; n26537
g26282 and n26450_not n26453_not ; n26538
g26283 and n26537 n26538 ; n26539
g26284 and n26537_not n26538_not ; n26540
g26285 and n26539_not n26540_not ; n26541
g26286 and b[62] n9339 ; n26542
g26287 and b[60] n9732 ; n26543
g26288 and b[61] n9334 ; n26544
g26289 and n26543_not n26544_not ; n26545
g26290 and n26542_not n26545 ; n26546
g26291 and n9342 n13370 ; n26547
g26292 and n26546 n26547_not ; n26548
g26293 and a[53] n26548_not ; n26549
g26294 and a[53] n26549_not ; n26550
g26295 and n26548_not n26549_not ; n26551
g26296 and n26550_not n26551_not ; n26552
g26297 and n26541 n26552_not ; n26553
g26298 and n26541 n26553_not ; n26554
g26299 and n26552_not n26553_not ; n26555
g26300 and n26554_not n26555_not ; n26556
g26301 and n26456_not n26460_not ; n26557
g26302 and b[63] n8715 ; n26558
g26303 and n8365_not n26558_not ; n26559
g26304 and n13797_not n26558_not ; n26560
g26305 and n26559_not n26560_not ; n26561
g26306 and a[50] n26561_not ; n26562
g26307 and a[50]_not n26561 ; n26563
g26308 and n26562_not n26563_not ; n26564
g26309 and n26557_not n26564_not ; n26565
g26310 and n26557 n26564 ; n26566
g26311 and n26565_not n26566_not ; n26567
g26312 and n26556_not n26567 ; n26568
g26313 and n26556_not n26568_not ; n26569
g26314 and n26567 n26568_not ; n26570
g26315 and n26569_not n26570_not ; n26571
g26316 and n26464_not n26467_not ; n26572
g26317 and n26571 n26572 ; n26573
g26318 and n26571_not n26572_not ; n26574
g26319 and n26573_not n26574_not ; n26575
g26320 and n26473_not n26476_not ; n26576
g26321 and n26575 n26576_not ; n26577
g26322 and n26575_not n26576 ; n26578
g26323 and n26577_not n26578_not ; f[113]
g26324 and n26531_not n26534_not ; n26580
g26325 and b[60] n10426 ; n26581
g26326 and b[58] n10796 ; n26582
g26327 and b[59] n10421 ; n26583
g26328 and n26582_not n26583_not ; n26584
g26329 and n26581_not n26584 ; n26585
g26330 and n10429 n12211 ; n26586
g26331 and n26585 n26586_not ; n26587
g26332 and a[56] n26587_not ; n26588
g26333 and a[56] n26588_not ; n26589
g26334 and n26587_not n26588_not ; n26590
g26335 and n26589_not n26590_not ; n26591
g26336 and n26515_not n26529_not ; n26592
g26337 and b[57] n11531 ; n26593
g26338 and b[55] n11896 ; n26594
g26339 and b[56] n11526 ; n26595
g26340 and n26594_not n26595_not ; n26596
g26341 and n26593_not n26596 ; n26597
g26342 and n11410 n11534 ; n26598
g26343 and n26597 n26598_not ; n26599
g26344 and a[59] n26599_not ; n26600
g26345 and a[59] n26600_not ; n26601
g26346 and n26599_not n26600_not ; n26602
g26347 and n26601_not n26602_not ; n26603
g26348 and b[54] n12668 ; n26604
g26349 and b[52] n13047 ; n26605
g26350 and b[53] n12663 ; n26606
g26351 and n26605_not n26606_not ; n26607
g26352 and n26604_not n26607 ; n26608
g26353 and n9998 n12671 ; n26609
g26354 and n26608 n26609_not ; n26610
g26355 and a[62] n26610_not ; n26611
g26356 and a[62] n26611_not ; n26612
g26357 and n26610_not n26611_not ; n26613
g26358 and n26612_not n26613_not ; n26614
g26359 and n26505_not n26509_not ; n26615
g26360 and b[50] n13903 ; n26616
g26361 and b[51] n13488_not ; n26617
g26362 and n26616_not n26617_not ; n26618
g26363 and a[50]_not n26618_not ; n26619
g26364 and a[50] n26618 ; n26620
g26365 and n26619_not n26620_not ; n26621
g26366 and n26422_not n26621 ; n26622
g26367 and n26422 n26621_not ; n26623
g26368 and n26622_not n26623_not ; n26624
g26369 and n26615_not n26624 ; n26625
g26370 and n26615_not n26625_not ; n26626
g26371 and n26624 n26625_not ; n26627
g26372 and n26626_not n26627_not ; n26628
g26373 and n26614_not n26628_not ; n26629
g26374 and n26614 n26627_not ; n26630
g26375 and n26626_not n26630 ; n26631
g26376 and n26629_not n26631_not ; n26632
g26377 and n26603_not n26632 ; n26633
g26378 and n26603_not n26633_not ; n26634
g26379 and n26632 n26633_not ; n26635
g26380 and n26634_not n26635_not ; n26636
g26381 and n26592_not n26636_not ; n26637
g26382 and n26592 n26635_not ; n26638
g26383 and n26634_not n26638 ; n26639
g26384 and n26637_not n26639_not ; n26640
g26385 and n26591_not n26640 ; n26641
g26386 and n26591 n26640_not ; n26642
g26387 and n26641_not n26642_not ; n26643
g26388 and n26580_not n26643 ; n26644
g26389 and n26580 n26643_not ; n26645
g26390 and n26644_not n26645_not ; n26646
g26391 and b[63] n9339 ; n26647
g26392 and b[61] n9732 ; n26648
g26393 and b[62] n9334 ; n26649
g26394 and n26648_not n26649_not ; n26650
g26395 and n26647_not n26650 ; n26651
g26396 and n9342 n13771 ; n26652
g26397 and n26651 n26652_not ; n26653
g26398 and a[53] n26653_not ; n26654
g26399 and a[53] n26654_not ; n26655
g26400 and n26653_not n26654_not ; n26656
g26401 and n26655_not n26656_not ; n26657
g26402 and n26646 n26657_not ; n26658
g26403 and n26646 n26658_not ; n26659
g26404 and n26657_not n26658_not ; n26660
g26405 and n26659_not n26660_not ; n26661
g26406 and n26540_not n26553_not ; n26662
g26407 and n26661 n26662 ; n26663
g26408 and n26661_not n26662_not ; n26664
g26409 and n26663_not n26664_not ; n26665
g26410 and n26565_not n26568_not ; n26666
g26411 and n26665_not n26666 ; n26667
g26412 and n26665 n26666_not ; n26668
g26413 and n26667_not n26668_not ; n26669
g26414 and n26574_not n26577_not ; n26670
g26415 and n26669 n26670_not ; n26671
g26416 and n26669_not n26670 ; n26672
g26417 and n26671_not n26672_not ; f[114]
g26418 and b[62] n9732 ; n26674
g26419 and b[63] n9334 ; n26675
g26420 and n26674_not n26675_not ; n26676
g26421 and n9342 n13800_not ; n26677
g26422 and n26676 n26677_not ; n26678
g26423 and a[53] n26678_not ; n26679
g26424 and a[53] n26679_not ; n26680
g26425 and n26678_not n26679_not ; n26681
g26426 and n26680_not n26681_not ; n26682
g26427 and n26641_not n26644_not ; n26683
g26428 and b[61] n10426 ; n26684
g26429 and b[59] n10796 ; n26685
g26430 and b[60] n10421 ; n26686
g26431 and n26685_not n26686_not ; n26687
g26432 and n26684_not n26687 ; n26688
g26433 and n10429 n12969 ; n26689
g26434 and n26688 n26689_not ; n26690
g26435 and a[56] n26690_not ; n26691
g26436 and a[56] n26691_not ; n26692
g26437 and n26690_not n26691_not ; n26693
g26438 and n26692_not n26693_not ; n26694
g26439 and n26633_not n26637_not ; n26695
g26440 and b[58] n11531 ; n26696
g26441 and b[56] n11896 ; n26697
g26442 and b[57] n11526 ; n26698
g26443 and n26697_not n26698_not ; n26699
g26444 and n26696_not n26699 ; n26700
g26445 and n11436 n11534 ; n26701
g26446 and n26700 n26701_not ; n26702
g26447 and a[59] n26702_not ; n26703
g26448 and a[59] n26703_not ; n26704
g26449 and n26702_not n26703_not ; n26705
g26450 and n26704_not n26705_not ; n26706
g26451 and n26625_not n26629_not ; n26707
g26452 and b[51] n13903 ; n26708
g26453 and b[52] n13488_not ; n26709
g26454 and n26708_not n26709_not ; n26710
g26455 and n26619_not n26622_not ; n26711
g26456 and n26710_not n26711 ; n26712
g26457 and n26710 n26711_not ; n26713
g26458 and n26712_not n26713_not ; n26714
g26459 and b[55] n12668 ; n26715
g26460 and b[53] n13047 ; n26716
g26461 and b[54] n12663 ; n26717
g26462 and n26716_not n26717_not ; n26718
g26463 and n26715_not n26718 ; n26719
g26464 and n10684 n12671 ; n26720
g26465 and n26719 n26720_not ; n26721
g26466 and a[62] n26721_not ; n26722
g26467 and a[62] n26722_not ; n26723
g26468 and n26721_not n26722_not ; n26724
g26469 and n26723_not n26724_not ; n26725
g26470 and n26714_not n26725 ; n26726
g26471 and n26714 n26725_not ; n26727
g26472 and n26726_not n26727_not ; n26728
g26473 and n26707_not n26728 ; n26729
g26474 and n26707 n26728_not ; n26730
g26475 and n26729_not n26730_not ; n26731
g26476 and n26706_not n26731 ; n26732
g26477 and n26706 n26731_not ; n26733
g26478 and n26732_not n26733_not ; n26734
g26479 and n26695_not n26734 ; n26735
g26480 and n26695_not n26735_not ; n26736
g26481 and n26734 n26735_not ; n26737
g26482 and n26736_not n26737_not ; n26738
g26483 and n26694_not n26738_not ; n26739
g26484 and n26694 n26737_not ; n26740
g26485 and n26736_not n26740 ; n26741
g26486 and n26739_not n26741_not ; n26742
g26487 and n26683_not n26742 ; n26743
g26488 and n26683 n26742_not ; n26744
g26489 and n26743_not n26744_not ; n26745
g26490 and n26682_not n26745 ; n26746
g26491 and n26745 n26746_not ; n26747
g26492 and n26682_not n26746_not ; n26748
g26493 and n26747_not n26748_not ; n26749
g26494 and n26658_not n26664_not ; n26750
g26495 and n26749 n26750 ; n26751
g26496 and n26749_not n26750_not ; n26752
g26497 and n26751_not n26752_not ; n26753
g26498 and n26668_not n26671_not ; n26754
g26499 and n26753 n26754_not ; n26755
g26500 and n26753_not n26754 ; n26756
g26501 and n26755_not n26756_not ; f[115]
g26502 and n26729_not n26732_not ; n26758
g26503 and n26713_not n26727_not ; n26759
g26504 and b[52] n13903 ; n26760
g26505 and b[53] n13488_not ; n26761
g26506 and n26760_not n26761_not ; n26762
g26507 and n26710 n26762_not ; n26763
g26508 and n26710_not n26762 ; n26764
g26509 and n26759_not n26764_not ; n26765
g26510 and n26763_not n26765 ; n26766
g26511 and n26759_not n26766_not ; n26767
g26512 and n26764_not n26766_not ; n26768
g26513 and n26763_not n26768 ; n26769
g26514 and n26767_not n26769_not ; n26770
g26515 and b[56] n12668 ; n26771
g26516 and b[54] n13047 ; n26772
g26517 and b[55] n12663 ; n26773
g26518 and n26772_not n26773_not ; n26774
g26519 and n26771_not n26774 ; n26775
g26520 and n10708 n12671 ; n26776
g26521 and n26775 n26776_not ; n26777
g26522 and a[62] n26777_not ; n26778
g26523 and a[62] n26778_not ; n26779
g26524 and n26777_not n26778_not ; n26780
g26525 and n26779_not n26780_not ; n26781
g26526 and n26770_not n26781 ; n26782
g26527 and n26770 n26781_not ; n26783
g26528 and n26782_not n26783_not ; n26784
g26529 and b[59] n11531 ; n26785
g26530 and b[57] n11896 ; n26786
g26531 and b[58] n11526 ; n26787
g26532 and n26786_not n26787_not ; n26788
g26533 and n26785_not n26788 ; n26789
g26534 and n11534 n12179 ; n26790
g26535 and n26789 n26790_not ; n26791
g26536 and a[59] n26791_not ; n26792
g26537 and a[59] n26792_not ; n26793
g26538 and n26791_not n26792_not ; n26794
g26539 and n26793_not n26794_not ; n26795
g26540 and n26784_not n26795_not ; n26796
g26541 and n26784 n26795 ; n26797
g26542 and n26796_not n26797_not ; n26798
g26543 and n26758 n26798_not ; n26799
g26544 and n26758_not n26798 ; n26800
g26545 and n26799_not n26800_not ; n26801
g26546 and b[62] n10426 ; n26802
g26547 and b[60] n10796 ; n26803
g26548 and b[61] n10421 ; n26804
g26549 and n26803_not n26804_not ; n26805
g26550 and n26802_not n26805 ; n26806
g26551 and n10429 n13370 ; n26807
g26552 and n26806 n26807_not ; n26808
g26553 and a[56] n26808_not ; n26809
g26554 and a[56] n26809_not ; n26810
g26555 and n26808_not n26809_not ; n26811
g26556 and n26810_not n26811_not ; n26812
g26557 and n26801 n26812_not ; n26813
g26558 and n26801 n26813_not ; n26814
g26559 and n26812_not n26813_not ; n26815
g26560 and n26814_not n26815_not ; n26816
g26561 and n26735_not n26739_not ; n26817
g26562 and b[63] n9732 ; n26818
g26563 and n9342_not n26818_not ; n26819
g26564 and n13797_not n26818_not ; n26820
g26565 and n26819_not n26820_not ; n26821
g26566 and a[53] n26821_not ; n26822
g26567 and a[53]_not n26821 ; n26823
g26568 and n26822_not n26823_not ; n26824
g26569 and n26817_not n26824_not ; n26825
g26570 and n26817 n26824 ; n26826
g26571 and n26825_not n26826_not ; n26827
g26572 and n26816_not n26827 ; n26828
g26573 and n26816_not n26828_not ; n26829
g26574 and n26827 n26828_not ; n26830
g26575 and n26829_not n26830_not ; n26831
g26576 and n26743_not n26746_not ; n26832
g26577 and n26831 n26832 ; n26833
g26578 and n26831_not n26832_not ; n26834
g26579 and n26833_not n26834_not ; n26835
g26580 and n26752_not n26755_not ; n26836
g26581 and n26835 n26836_not ; n26837
g26582 and n26835_not n26836 ; n26838
g26583 and n26837_not n26838_not ; f[116]
g26584 and n26834_not n26837_not ; n26840
g26585 and n26825_not n26828_not ; n26841
g26586 and n26800_not n26813_not ; n26842
g26587 and b[63] n10426 ; n26843
g26588 and b[61] n10796 ; n26844
g26589 and b[62] n10421 ; n26845
g26590 and n26844_not n26845_not ; n26846
g26591 and n26843_not n26846 ; n26847
g26592 and n10429 n13771 ; n26848
g26593 and n26847 n26848_not ; n26849
g26594 and a[56] n26849_not ; n26850
g26595 and a[56] n26850_not ; n26851
g26596 and n26849_not n26850_not ; n26852
g26597 and n26851_not n26852_not ; n26853
g26598 and n26842_not n26853_not ; n26854
g26599 and n26842_not n26854_not ; n26855
g26600 and n26853_not n26854_not ; n26856
g26601 and n26855_not n26856_not ; n26857
g26602 and n26770_not n26781_not ; n26858
g26603 and n26796_not n26858_not ; n26859
g26604 and b[60] n11531 ; n26860
g26605 and b[58] n11896 ; n26861
g26606 and b[59] n11526 ; n26862
g26607 and n26861_not n26862_not ; n26863
g26608 and n26860_not n26863 ; n26864
g26609 and n11534 n12211 ; n26865
g26610 and n26864 n26865_not ; n26866
g26611 and a[59] n26866_not ; n26867
g26612 and a[59] n26867_not ; n26868
g26613 and n26866_not n26867_not ; n26869
g26614 and n26868_not n26869_not ; n26870
g26615 and a[53] n26762_not ; n26871
g26616 and a[53]_not n26762 ; n26872
g26617 and n26871_not n26872_not ; n26873
g26618 and b[53] n13903 ; n26874
g26619 and b[54] n13488_not ; n26875
g26620 and n26874_not n26875_not ; n26876
g26621 and n26873 n26876 ; n26877
g26622 and n26873_not n26876_not ; n26878
g26623 and n26877_not n26878_not ; n26879
g26624 and b[57] n12668 ; n26880
g26625 and b[55] n13047 ; n26881
g26626 and b[56] n12663 ; n26882
g26627 and n26881_not n26882_not ; n26883
g26628 and n26880_not n26883 ; n26884
g26629 and n11410 n12671 ; n26885
g26630 and n26884 n26885_not ; n26886
g26631 and a[62] n26886_not ; n26887
g26632 and a[62] n26887_not ; n26888
g26633 and n26886_not n26887_not ; n26889
g26634 and n26888_not n26889_not ; n26890
g26635 and n26879 n26890_not ; n26891
g26636 and n26879 n26891_not ; n26892
g26637 and n26890_not n26891_not ; n26893
g26638 and n26892_not n26893_not ; n26894
g26639 and n26768_not n26894_not ; n26895
g26640 and n26768 n26894 ; n26896
g26641 and n26895_not n26896_not ; n26897
g26642 and n26870_not n26897 ; n26898
g26643 and n26870_not n26898_not ; n26899
g26644 and n26897 n26898_not ; n26900
g26645 and n26899_not n26900_not ; n26901
g26646 and n26859_not n26901_not ; n26902
g26647 and n26859_not n26902_not ; n26903
g26648 and n26901_not n26902_not ; n26904
g26649 and n26903_not n26904_not ; n26905
g26650 and n26857_not n26905 ; n26906
g26651 and n26857 n26905_not ; n26907
g26652 and n26906_not n26907_not ; n26908
g26653 and n26841_not n26908_not ; n26909
g26654 and n26841 n26908 ; n26910
g26655 and n26909_not n26910_not ; n26911
g26656 and n26840_not n26911 ; n26912
g26657 and n26840 n26911_not ; n26913
g26658 and n26912_not n26913_not ; f[117]
g26659 and b[62] n10796 ; n26915
g26660 and b[63] n10421 ; n26916
g26661 and n26915_not n26916_not ; n26917
g26662 and n10429 n13800_not ; n26918
g26663 and n26917 n26918_not ; n26919
g26664 and a[56] n26919_not ; n26920
g26665 and a[56] n26920_not ; n26921
g26666 and n26919_not n26920_not ; n26922
g26667 and n26921_not n26922_not ; n26923
g26668 and n26898_not n26902_not ; n26924
g26669 and b[61] n11531 ; n26925
g26670 and b[59] n11896 ; n26926
g26671 and b[60] n11526 ; n26927
g26672 and n26926_not n26927_not ; n26928
g26673 and n26925_not n26928 ; n26929
g26674 and n11534 n12969 ; n26930
g26675 and n26929 n26930_not ; n26931
g26676 and a[59] n26931_not ; n26932
g26677 and a[59] n26932_not ; n26933
g26678 and n26931_not n26932_not ; n26934
g26679 and n26933_not n26934_not ; n26935
g26680 and n26891_not n26895_not ; n26936
g26681 and b[54] n13903 ; n26937
g26682 and b[55] n13488_not ; n26938
g26683 and n26937_not n26938_not ; n26939
g26684 and a[53]_not n26762_not ; n26940
g26685 and n26878_not n26940_not ; n26941
g26686 and n26939 n26941_not ; n26942
g26687 and n26939_not n26941 ; n26943
g26688 and n26942_not n26943_not ; n26944
g26689 and b[58] n12668 ; n26945
g26690 and b[56] n13047 ; n26946
g26691 and b[57] n12663 ; n26947
g26692 and n26946_not n26947_not ; n26948
g26693 and n26945_not n26948 ; n26949
g26694 and n12671_not n26949 ; n26950
g26695 and n11436_not n26949 ; n26951
g26696 and n26950_not n26951_not ; n26952
g26697 and a[62] n26952_not ; n26953
g26698 and a[62]_not n26952 ; n26954
g26699 and n26953_not n26954_not ; n26955
g26700 and n26944 n26955_not ; n26956
g26701 and n26944_not n26955 ; n26957
g26702 and n26956_not n26957_not ; n26958
g26703 and n26936_not n26958 ; n26959
g26704 and n26936_not n26959_not ; n26960
g26705 and n26958 n26959_not ; n26961
g26706 and n26960_not n26961_not ; n26962
g26707 and n26935_not n26962_not ; n26963
g26708 and n26935 n26961_not ; n26964
g26709 and n26960_not n26964 ; n26965
g26710 and n26963_not n26965_not ; n26966
g26711 and n26924_not n26966 ; n26967
g26712 and n26924 n26966_not ; n26968
g26713 and n26967_not n26968_not ; n26969
g26714 and n26923_not n26969 ; n26970
g26715 and n26969 n26970_not ; n26971
g26716 and n26923_not n26970_not ; n26972
g26717 and n26971_not n26972_not ; n26973
g26718 and n26857_not n26905_not ; n26974
g26719 and n26854_not n26974_not ; n26975
g26720 and n26973_not n26975_not ; n26976
g26721 and n26973_not n26976_not ; n26977
g26722 and n26975_not n26976_not ; n26978
g26723 and n26977_not n26978_not ; n26979
g26724 and n26909_not n26912_not ; n26980
g26725 and n26979_not n26980_not ; n26981
g26726 and n26979 n26980 ; n26982
g26727 and n26981_not n26982_not ; f[118]
g26728 and b[59] n12668 ; n26984
g26729 and b[57] n13047 ; n26985
g26730 and b[58] n12663 ; n26986
g26731 and n26985_not n26986_not ; n26987
g26732 and n26984_not n26987 ; n26988
g26733 and n12179 n12671 ; n26989
g26734 and n26988 n26989_not ; n26990
g26735 and a[62] n26990_not ; n26991
g26736 and a[62] n26991_not ; n26992
g26737 and n26990_not n26991_not ; n26993
g26738 and n26992_not n26993_not ; n26994
g26739 and b[55] n13903 ; n26995
g26740 and b[56] n13488_not ; n26996
g26741 and n26995_not n26996_not ; n26997
g26742 and n26939 n26997_not ; n26998
g26743 and n26939 n26998_not ; n26999
g26744 and n26997_not n26998_not ; n27000
g26745 and n26999_not n27000_not ; n27001
g26746 and n26994_not n27001_not ; n27002
g26747 and n26994_not n27002_not ; n27003
g26748 and n27001_not n27002_not ; n27004
g26749 and n27003_not n27004_not ; n27005
g26750 and n26942_not n26956_not ; n27006
g26751 and n27005 n27006 ; n27007
g26752 and n27005_not n27006_not ; n27008
g26753 and n27007_not n27008_not ; n27009
g26754 and b[62] n11531 ; n27010
g26755 and b[60] n11896 ; n27011
g26756 and b[61] n11526 ; n27012
g26757 and n27011_not n27012_not ; n27013
g26758 and n27010_not n27013 ; n27014
g26759 and n11534 n13370 ; n27015
g26760 and n27014 n27015_not ; n27016
g26761 and a[59] n27016_not ; n27017
g26762 and a[59] n27017_not ; n27018
g26763 and n27016_not n27017_not ; n27019
g26764 and n27018_not n27019_not ; n27020
g26765 and n27009 n27020_not ; n27021
g26766 and n27009 n27021_not ; n27022
g26767 and n27020_not n27021_not ; n27023
g26768 and n27022_not n27023_not ; n27024
g26769 and n26959_not n26963_not ; n27025
g26770 and b[63] n10796 ; n27026
g26771 and n10429_not n27026_not ; n27027
g26772 and n13797_not n27026_not ; n27028
g26773 and n27027_not n27028_not ; n27029
g26774 and a[56] n27029_not ; n27030
g26775 and a[56]_not n27029 ; n27031
g26776 and n27030_not n27031_not ; n27032
g26777 and n27025_not n27032_not ; n27033
g26778 and n27025 n27032 ; n27034
g26779 and n27033_not n27034_not ; n27035
g26780 and n27024_not n27035 ; n27036
g26781 and n27024_not n27036_not ; n27037
g26782 and n27035 n27036_not ; n27038
g26783 and n27037_not n27038_not ; n27039
g26784 and n26967_not n26970_not ; n27040
g26785 and n27039 n27040 ; n27041
g26786 and n27039_not n27040_not ; n27042
g26787 and n27041_not n27042_not ; n27043
g26788 and n26976_not n26981_not ; n27044
g26789 and n27043 n27044_not ; n27045
g26790 and n27043_not n27044 ; n27046
g26791 and n27045_not n27046_not ; f[119]
g26792 and n27008_not n27021_not ; n27048
g26793 and b[63] n11531 ; n27049
g26794 and b[61] n11896 ; n27050
g26795 and b[62] n11526 ; n27051
g26796 and n27050_not n27051_not ; n27052
g26797 and n27049_not n27052 ; n27053
g26798 and n11534 n13771 ; n27054
g26799 and n27053 n27054_not ; n27055
g26800 and a[59] n27055_not ; n27056
g26801 and a[59] n27056_not ; n27057
g26802 and n27055_not n27056_not ; n27058
g26803 and n27057_not n27058_not ; n27059
g26804 and n27048_not n27059_not ; n27060
g26805 and n27048_not n27060_not ; n27061
g26806 and n27059_not n27060_not ; n27062
g26807 and n27061_not n27062_not ; n27063
g26808 and b[56] n13903 ; n27064
g26809 and b[57] n13488_not ; n27065
g26810 and n27064_not n27065_not ; n27066
g26811 and a[56]_not n27066_not ; n27067
g26812 and a[56]_not n27067_not ; n27068
g26813 and n27066_not n27067_not ; n27069
g26814 and n27068_not n27069_not ; n27070
g26815 and n26939_not n27070_not ; n27071
g26816 and n26939_not n27071_not ; n27072
g26817 and n27070_not n27071_not ; n27073
g26818 and n27072_not n27073_not ; n27074
g26819 and n26998_not n27002_not ; n27075
g26820 and n27074 n27075 ; n27076
g26821 and n27074_not n27075_not ; n27077
g26822 and n27076_not n27077_not ; n27078
g26823 and b[60] n12668 ; n27079
g26824 and b[58] n13047 ; n27080
g26825 and b[59] n12663 ; n27081
g26826 and n27080_not n27081_not ; n27082
g26827 and n27079_not n27082 ; n27083
g26828 and n12211 n12671 ; n27084
g26829 and n27083 n27084_not ; n27085
g26830 and a[62] n27085_not ; n27086
g26831 and a[62] n27086_not ; n27087
g26832 and n27085_not n27086_not ; n27088
g26833 and n27087_not n27088_not ; n27089
g26834 and n27078 n27089_not ; n27090
g26835 and n27078_not n27089 ; n27091
g26836 and n27063_not n27091_not ; n27092
g26837 and n27090_not n27092 ; n27093
g26838 and n27063_not n27093_not ; n27094
g26839 and n27091_not n27093_not ; n27095
g26840 and n27090_not n27095 ; n27096
g26841 and n27094_not n27096_not ; n27097
g26842 and n27033_not n27036_not ; n27098
g26843 and n27097 n27098 ; n27099
g26844 and n27097_not n27098_not ; n27100
g26845 and n27099_not n27100_not ; n27101
g26846 and n27042_not n27045_not ; n27102
g26847 and n27101 n27102_not ; n27103
g26848 and n27101_not n27102 ; n27104
g26849 and n27103_not n27104_not ; f[120]
g26850 and n27077_not n27090_not ; n27106
g26851 and b[57] n13903 ; n27107
g26852 and b[58] n13488_not ; n27108
g26853 and n27107_not n27108_not ; n27109
g26854 and n27067_not n27071_not ; n27110
g26855 and n27109_not n27110 ; n27111
g26856 and n27109 n27110_not ; n27112
g26857 and n27111_not n27112_not ; n27113
g26858 and b[61] n12668 ; n27114
g26859 and b[59] n13047 ; n27115
g26860 and b[60] n12663 ; n27116
g26861 and n27115_not n27116_not ; n27117
g26862 and n27114_not n27117 ; n27118
g26863 and n12671_not n27118 ; n27119
g26864 and n12969_not n27118 ; n27120
g26865 and n27119_not n27120_not ; n27121
g26866 and a[62] n27121_not ; n27122
g26867 and a[62]_not n27121 ; n27123
g26868 and n27122_not n27123_not ; n27124
g26869 and n27113 n27124_not ; n27125
g26870 and n27113_not n27124 ; n27126
g26871 and n27125_not n27126_not ; n27127
g26872 and n27106_not n27127 ; n27128
g26873 and n27106 n27127_not ; n27129
g26874 and n27128_not n27129_not ; n27130
g26875 and b[62] n11896 ; n27131
g26876 and b[63] n11526 ; n27132
g26877 and n27131_not n27132_not ; n27133
g26878 and n11534 n13800_not ; n27134
g26879 and n27133 n27134_not ; n27135
g26880 and a[59] n27135_not ; n27136
g26881 and a[59] n27136_not ; n27137
g26882 and n27135_not n27136_not ; n27138
g26883 and n27137_not n27138_not ; n27139
g26884 and n27130 n27139_not ; n27140
g26885 and n27130 n27140_not ; n27141
g26886 and n27139_not n27140_not ; n27142
g26887 and n27141_not n27142_not ; n27143
g26888 and n27060_not n27093_not ; n27144
g26889 and n27143 n27144 ; n27145
g26890 and n27143_not n27144_not ; n27146
g26891 and n27145_not n27146_not ; n27147
g26892 and n27100_not n27103_not ; n27148
g26893 and n27147 n27148_not ; n27149
g26894 and n27147_not n27148 ; n27150
g26895 and n27149_not n27150_not ; f[121]
g26896 and n27146_not n27149_not ; n27152
g26897 and n27128_not n27140_not ; n27153
g26898 and n27112_not n27125_not ; n27154
g26899 and b[58] n13903 ; n27155
g26900 and b[59] n13488_not ; n27156
g26901 and n27155_not n27156_not ; n27157
g26902 and n27109 n27157_not ; n27158
g26903 and n27109_not n27157 ; n27159
g26904 and n27154_not n27159_not ; n27160
g26905 and n27158_not n27160 ; n27161
g26906 and n27154_not n27161_not ; n27162
g26907 and n27159_not n27161_not ; n27163
g26908 and n27158_not n27163 ; n27164
g26909 and n27162_not n27164_not ; n27165
g26910 and b[62] n12668 ; n27166
g26911 and b[60] n13047 ; n27167
g26912 and b[61] n12663 ; n27168
g26913 and n27167_not n27168_not ; n27169
g26914 and n27166_not n27169 ; n27170
g26915 and n12671 n13370 ; n27171
g26916 and n27170 n27171_not ; n27172
g26917 and a[62] n27172_not ; n27173
g26918 and a[62] n27173_not ; n27174
g26919 and n27172_not n27173_not ; n27175
g26920 and n27174_not n27175_not ; n27176
g26921 and b[63] n11896 ; n27177
g26922 and n11534 n13797 ; n27178
g26923 and n27177_not n27178_not ; n27179
g26924 and a[59] n27179_not ; n27180
g26925 and a[59] n27180_not ; n27181
g26926 and n27179_not n27180_not ; n27182
g26927 and n27181_not n27182_not ; n27183
g26928 and n27176_not n27183_not ; n27184
g26929 and n27176_not n27184_not ; n27185
g26930 and n27183_not n27184_not ; n27186
g26931 and n27185_not n27186_not ; n27187
g26932 and n27165_not n27187 ; n27188
g26933 and n27165 n27187_not ; n27189
g26934 and n27188_not n27189_not ; n27190
g26935 and n27153_not n27190_not ; n27191
g26936 and n27153_not n27191_not ; n27192
g26937 and n27190_not n27191_not ; n27193
g26938 and n27192_not n27193_not ; n27194
g26939 and n27152_not n27194_not ; n27195
g26940 and n27152 n27193_not ; n27196
g26941 and n27192_not n27196 ; n27197
g26942 and n27195_not n27197_not ; f[122]
g26943 and n27191_not n27195_not ; n27199
g26944 and n27165_not n27187_not ; n27200
g26945 and n27184_not n27200_not ; n27201
g26946 and a[59] n27157_not ; n27202
g26947 and a[59]_not n27157 ; n27203
g26948 and n27202_not n27203_not ; n27204
g26949 and b[59] n13903 ; n27205
g26950 and b[60] n13488_not ; n27206
g26951 and n27205_not n27206_not ; n27207
g26952 and n27204 n27207 ; n27208
g26953 and n27204_not n27207_not ; n27209
g26954 and n27208_not n27209_not ; n27210
g26955 and b[63] n12668 ; n27211
g26956 and b[61] n13047 ; n27212
g26957 and b[62] n12663 ; n27213
g26958 and n27212_not n27213_not ; n27214
g26959 and n27211_not n27214 ; n27215
g26960 and n12671 n13771 ; n27216
g26961 and n27215 n27216_not ; n27217
g26962 and a[62] n27217_not ; n27218
g26963 and a[62] n27218_not ; n27219
g26964 and n27217_not n27218_not ; n27220
g26965 and n27219_not n27220_not ; n27221
g26966 and n27210 n27221_not ; n27222
g26967 and n27210 n27222_not ; n27223
g26968 and n27221_not n27222_not ; n27224
g26969 and n27223_not n27224_not ; n27225
g26970 and n27163_not n27225_not ; n27226
g26971 and n27163 n27225 ; n27227
g26972 and n27226_not n27227_not ; n27228
g26973 and n27201_not n27228 ; n27229
g26974 and n27201_not n27229_not ; n27230
g26975 and n27228 n27229_not ; n27231
g26976 and n27230_not n27231_not ; n27232
g26977 and n27199_not n27232_not ; n27233
g26978 and n27199 n27231_not ; n27234
g26979 and n27230_not n27234 ; n27235
g26980 and n27233_not n27235_not ; f[123]
g26981 and n27229_not n27233_not ; n27237
g26982 and n27222_not n27226_not ; n27238
g26983 and b[60] n13903 ; n27239
g26984 and b[61] n13488_not ; n27240
g26985 and n27239_not n27240_not ; n27241
g26986 and a[59]_not n27157_not ; n27242
g26987 and n27209_not n27242_not ; n27243
g26988 and n27241 n27243_not ; n27244
g26989 and n27241_not n27243 ; n27245
g26990 and n27244_not n27245_not ; n27246
g26991 and b[62] n13047 ; n27247
g26992 and b[63] n12663 ; n27248
g26993 and n27247_not n27248_not ; n27249
g26994 and n12671_not n27249 ; n27250
g26995 and n13800 n27249 ; n27251
g26996 and n27250_not n27251_not ; n27252
g26997 and a[62] n27252_not ; n27253
g26998 and a[62]_not n27252 ; n27254
g26999 and n27253_not n27254_not ; n27255
g27000 and n27246 n27255_not ; n27256
g27001 and n27246_not n27255 ; n27257
g27002 and n27256_not n27257_not ; n27258
g27003 and n27238_not n27258 ; n27259
g27004 and n27238_not n27259_not ; n27260
g27005 and n27258 n27259_not ; n27261
g27006 and n27260_not n27261_not ; n27262
g27007 and n27237_not n27262_not ; n27263
g27008 and n27237 n27261_not ; n27264
g27009 and n27260_not n27264 ; n27265
g27010 and n27263_not n27265_not ; f[124]
g27011 and n27259_not n27263_not ; n27267
g27012 and n27244_not n27256_not ; n27268
g27013 and b[61] n13903 ; n27269
g27014 and b[62] n13488_not ; n27270
g27015 and n27269_not n27270_not ; n27271
g27016 and n27241 n27271_not ; n27272
g27017 and n27241_not n27271 ; n27273
g27018 and n27272_not n27273_not ; n27274
g27019 and b[63] n13047 ; n27275
g27020 and n12671_not n27275_not ; n27276
g27021 and n13797_not n27275_not ; n27277
g27022 and n27276_not n27277_not ; n27278
g27023 and a[62] n27278_not ; n27279
g27024 and a[62]_not n27278 ; n27280
g27025 and n27279_not n27280_not ; n27281
g27026 and n27274 n27281_not ; n27282
g27027 and n27274_not n27281 ; n27283
g27028 and n27282_not n27283_not ; n27284
g27029 and n27268_not n27284 ; n27285
g27030 and n27268_not n27285_not ; n27286
g27031 and n27284 n27285_not ; n27287
g27032 and n27286_not n27287_not ; n27288
g27033 and n27267_not n27288_not ; n27289
g27034 and n27267 n27287_not ; n27290
g27035 and n27286_not n27290 ; n27291
g27036 and n27289_not n27291_not ; f[125]
g27037 and n27285_not n27289_not ; n27293
g27038 and n27272_not n27282_not ; n27294
g27039 and b[62] n13903 ; n27295
g27040 and b[63] n13488_not ; n27296
g27041 and n27295_not n27296_not ; n27297
g27042 and a[62]_not n27297_not ; n27298
g27043 and a[62] n27297 ; n27299
g27044 and n27298_not n27299_not ; n27300
g27045 and n27241_not n27300 ; n27301
g27046 and n27241 n27300_not ; n27302
g27047 and n27301_not n27302_not ; n27303
g27048 and n27294_not n27303 ; n27304
g27049 and n27294 n27303_not ; n27305
g27050 and n27304_not n27305_not ; n27306
g27051 and n27293_not n27306 ; n27307
g27052 and n27293 n27306_not ; n27308
g27053 and n27307_not n27308_not ; f[126]
g27054 and n27298_not n27301_not ; n27310
g27055 and b[63] n13903 ; n27311
g27056 and n27310_not n27311 ; n27312
g27057 and n27310 n27311_not ; n27313
g27058 and n27312_not n27313_not ; n27314
g27059 and n27304_not n27307_not ; n27315
g27060 and n27314 n27315 ; n27316
g27061 and n27314_not n27315_not ; n27317
g27062 and n27316_not n27317_not ; f[127]
g27063 not n300 ; n300_not
g27064 not n301 ; n301_not
g27065 not n400 ; n400_not
g27066 not n401 ; n401_not
g27067 not n302 ; n302_not
g27068 not n311 ; n311_not
g27069 not n320 ; n320_not
g27070 not n500 ; n500_not
g27071 not n410 ; n410_not
g27072 not n321 ; n321_not
g27073 not n600 ; n600_not
g27074 not n330 ; n330_not
g27075 not n312 ; n312_not
g27076 not n303 ; n303_not
g27077 not n420 ; n420_not
g27078 not n501 ; n501_not
g27079 not n411 ; n411_not
g27080 not n510 ; n510_not
g27081 not n313 ; n313_not
g27082 not n331 ; n331_not
g27083 not n421 ; n421_not
g27084 not n610 ; n610_not
g27085 not n340 ; n340_not
g27086 not n502 ; n502_not
g27087 not n430 ; n430_not
g27088 not n304 ; n304_not
g27089 not n412 ; n412_not
g27090 not n601 ; n601_not
g27091 not n520 ; n520_not
g27092 not n322 ; n322_not
g27093 not n332 ; n332_not
g27094 not n314 ; n314_not
g27095 not n440 ; n440_not
g27096 not n530 ; n530_not
g27097 not n620 ; n620_not
g27098 not n710 ; n710_not
g27099 not n323 ; n323_not
g27100 not n503 ; n503_not
g27101 not n431 ; n431_not
g27102 not n404 ; n404_not
g27103 not n611 ; n611_not
g27104 not n512 ; n512_not
g27105 not n422 ; n422_not
g27106 not n341 ; n341_not
g27107 not n413 ; n413_not
g27108 not n521 ; n521_not
g27109 not n800 ; n800_not
g27110 not n602 ; n602_not
g27111 not n701 ; n701_not
g27112 not n350 ; n350_not
g27113 not n522 ; n522_not
g27114 not n324 ; n324_not
g27115 not n630 ; n630_not
g27116 not n720 ; n720_not
g27117 not n450 ; n450_not
g27118 not n342 ; n342_not
g27119 not n333 ; n333_not
g27120 not n414 ; n414_not
g27121 not n351 ; n351_not
g27122 not n405 ; n405_not
g27123 not n900 ; n900_not
g27124 not n360 ; n360_not
g27125 not n423 ; n423_not
g27126 not n441 ; n441_not
g27127 not n711 ; n711_not
g27128 not n306 ; n306_not
g27129 not n504 ; n504_not
g27130 not n270 ; n270_not
g27131 not n531 ; n531_not
g27132 not n315 ; n315_not
g27133 not n432 ; n432_not
g27134 not n612 ; n612_not
g27135 not n801 ; n801_not
g27136 not n505 ; n505_not
g27137 not n361 ; n361_not
g27138 not n712 ; n712_not
g27139 not n514 ; n514_not
g27140 not n352 ; n352_not
g27141 not n703 ; n703_not
g27142 not n640 ; n640_not
g27143 not n370 ; n370_not
g27144 not n802 ; n802_not
g27145 not n901 ; n901_not
g27146 not n613 ; n613_not
g27147 not n460 ; n460_not
g27148 not n433 ; n433_not
g27149 not n262 ; n262_not
g27150 not n442 ; n442_not
g27151 not n271 ; n271_not
g27152 not n550 ; n550_not
g27153 not n280 ; n280_not
g27154 not n721 ; n721_not
g27155 not n343 ; n343_not
g27156 not n316 ; n316_not
g27157 not n415 ; n415_not
g27158 not n325 ; n325_not
g27159 not n820 ; n820_not
g27160 not n307 ; n307_not
g27161 not n532 ; n532_not
g27162 not n910 ; n910_not
g27163 not n632 ; n632_not
g27164 not n803 ; n803_not
g27165 not n533 ; n533_not
g27166 not n272 ; n272_not
g27167 not n614 ; n614_not
g27168 not n461 ; n461_not
g27169 not n623 ; n623_not
g27170 not n443 ; n443_not
g27171 not n434 ; n434_not
g27172 not n821 ; n821_not
g27173 not n425 ; n425_not
g27174 not n380 ; n380_not
g27175 not n470 ; n470_not
g27176 not n812 ; n812_not
g27177 not n605 ; n605_not
g27178 not n722 ; n722_not
g27179 not n524 ; n524_not
g27180 not n326 ; n326_not
g27181 not n317 ; n317_not
g27182 not n290 ; n290_not
g27183 not n308 ; n308_not
g27184 not n911 ; n911_not
g27185 not n542 ; n542_not
g27186 not n704 ; n704_not
g27187 not n902 ; n902_not
g27188 not n551 ; n551_not
g27189 not n560 ; n560_not
g27190 not n263 ; n263_not
g27191 not n344 ; n344_not
g27192 not n641 ; n641_not
g27193 not n740 ; n740_not
g27194 not n353 ; n353_not
g27195 not n371 ; n371_not
g27196 not n713 ; n713_not
g27197 not n920 ; n920_not
g27198 not n515 ; n515_not
g27199 not n335 ; n335_not
g27200 not n650 ; n650_not
g27201 not n813 ; n813_not
g27202 not n462 ; n462_not
g27203 not n606 ; n606_not
g27204 not n732 ; n732_not
g27205 not n525 ; n525_not
g27206 not n561 ; n561_not
g27207 not n453 ; n453_not
g27208 not n714 ; n714_not
g27209 not n444 ; n444_not
g27210 not n741 ; n741_not
g27211 not n552 ; n552_not
g27212 not n507 ; n507_not
g27213 not n804 ; n804_not
g27214 not n480 ; n480_not
g27215 not n534 ; n534_not
g27216 not n570 ; n570_not
g27217 not n822 ; n822_not
g27218 not n516 ; n516_not
g27219 not n543 ; n543_not
g27220 not n417 ; n417_not
g27221 not n282 ; n282_not
g27222 not n372 ; n372_not
g27223 not n291 ; n291_not
g27224 not n705 ; n705_not
g27225 not n408 ; n408_not
g27226 not n831 ; n831_not
g27227 not n840 ; n840_not
g27228 not n660 ; n660_not
g27229 not n912 ; n912_not
g27230 not n390 ; n390_not
g27231 not n633 ; n633_not
g27232 not n327 ; n327_not
g27233 not n381 ; n381_not
g27234 not n336 ; n336_not
g27235 not n642 ; n642_not
g27236 not n345 ; n345_not
g27237 not n363 ; n363_not
g27238 not n354 ; n354_not
g27239 not n930 ; n930_not
g27240 not n615 ; n615_not
g27241 not n723 ; n723_not
g27242 not n264 ; n264_not
g27243 not n435 ; n435_not
g27244 not n624 ; n624_not
g27245 not n426 ; n426_not
g27246 not n273 ; n273_not
g27247 not n903 ; n903_not
g27248 not n328 ; n328_not
g27249 not n292 ; n292_not
g27250 not n337 ; n337_not
g27251 not n265 ; n265_not
g27252 not n661 ; n661_not
g27253 not n652 ; n652_not
g27254 not n913 ; n913_not
g27255 not n742 ; n742_not
g27256 not n562 ; n562_not
g27257 not n571 ; n571_not
g27258 not n760 ; n760_not
g27259 not n517 ; n517_not
g27260 not n526 ; n526_not
g27261 not n319 ; n319_not
g27262 not n580 ; n580_not
g27263 not n904 ; n904_not
g27264 not n274 ; n274_not
g27265 not n940 ; n940_not
g27266 not n706 ; n706_not
g27267 not n490 ; n490_not
g27268 not n553 ; n553_not
g27269 not n472 ; n472_not
g27270 not n535 ; n535_not
g27271 not n814 ; n814_not
g27272 not n805 ; n805_not
g27273 not n409 ; n409_not
g27274 not n481 ; n481_not
g27275 not n931 ; n931_not
g27276 not n625 ; n625_not
g27277 not n607 ; n607_not
g27278 not n418 ; n418_not
g27279 not n724 ; n724_not
g27280 not n832 ; n832_not
g27281 not n427 ; n427_not
g27282 not n436 ; n436_not
g27283 not n751 ; n751_not
g27284 not n463 ; n463_not
g27285 not n445 ; n445_not
g27286 not n616 ; n616_not
g27287 not n823 ; n823_not
g27288 not n454 ; n454_not
g27289 not n373 ; n373_not
g27290 not n508 ; n508_not
g27291 not n634 ; n634_not
g27292 not n850 ; n850_not
g27293 not n715 ; n715_not
g27294 not n733 ; n733_not
g27295 not n355 ; n355_not
g27296 not n391 ; n391_not
g27297 not n841 ; n841_not
g27298 not n950 ; n950_not
g27299 not n680 ; n680_not
g27300 not n941 ; n941_not
g27301 not n743 ; n743_not
g27302 not n716 ; n716_not
g27303 not n581 ; n581_not
g27304 not n653 ; n653_not
g27305 not n590 ; n590_not
g27306 not n761 ; n761_not
g27307 not n608 ; n608_not
g27308 not n635 ; n635_not
g27309 not n662 ; n662_not
g27310 not n572 ; n572_not
g27311 not n734 ; n734_not
g27312 not n725 ; n725_not
g27313 not n707 ; n707_not
g27314 not n482 ; n482_not
g27315 not n626 ; n626_not
g27316 not n365 ; n365_not
g27317 not n617 ; n617_not
g27318 not n536 ; n536_not
g27319 not n329 ; n329_not
g27320 not n347 ; n347_not
g27321 not n752 ; n752_not
g27322 not n491 ; n491_not
g27323 not n356 ; n356_not
g27324 not n923 ; n923_not
g27325 not n815 ; n815_not
g27326 not n455 ; n455_not
g27327 not n473 ; n473_not
g27328 not n464 ; n464_not
g27329 not n806 ; n806_not
g27330 not n824 ; n824_not
g27331 not n392 ; n392_not
g27332 not n860 ; n860_not
g27333 not n851 ; n851_not
g27334 not n446 ; n446_not
g27335 not n428 ; n428_not
g27336 not n419 ; n419_not
g27337 not n833 ; n833_not
g27338 not n383 ; n383_not
g27339 not n932 ; n932_not
g27340 not n275 ; n275_not
g27341 not n527 ; n527_not
g27342 not n905 ; n905_not
g27343 not n257 ; n257_not
g27344 not n518 ; n518_not
g27345 not n563 ; n563_not
g27346 not n509 ; n509_not
g27347 not n914 ; n914_not
g27348 not n276 ; n276_not
g27349 not n636 ; n636_not
g27350 not n663 ; n663_not
g27351 not n681 ; n681_not
g27352 not n267 ; n267_not
g27353 not n672 ; n672_not
g27354 not n960 ; n960_not
g27355 not n942 ; n942_not
g27356 not n384 ; n384_not
g27357 not n843 ; n843_not
g27358 not n258 ; n258_not
g27359 not n708 ; n708_not
g27360 not n654 ; n654_not
g27361 not n348 ; n348_not
g27362 not n366 ; n366_not
g27363 not n645 ; n645_not
g27364 not n690 ; n690_not
g27365 not n294 ; n294_not
g27366 not n285 ; n285_not
g27367 not n924 ; n924_not
g27368 not n375 ; n375_not
g27369 not n717 ; n717_not
g27370 not n861 ; n861_not
g27371 not n816 ; n816_not
g27372 not n483 ; n483_not
g27373 not n807 ; n807_not
g27374 not n492 ; n492_not
g27375 not n429 ; n429_not
g27376 not n591 ; n591_not
g27377 not n735 ; n735_not
g27378 not n519 ; n519_not
g27379 not n726 ; n726_not
g27380 not n582 ; n582_not
g27381 not n744 ; n744_not
g27382 not n528 ; n528_not
g27383 not n537 ; n537_not
g27384 not n546 ; n546_not
g27385 not n753 ; n753_not
g27386 not n555 ; n555_not
g27387 not n564 ; n564_not
g27388 not n762 ; n762_not
g27389 not n618 ; n618_not
g27390 not n627 ; n627_not
g27391 not n825 ; n825_not
g27392 not n456 ; n456_not
g27393 not n447 ; n447_not
g27394 not n465 ; n465_not
g27395 not n393 ; n393_not
g27396 not n474 ; n474_not
g27397 not n933 ; n933_not
g27398 not n609 ; n609_not
g27399 not n745 ; n745_not
g27400 not n682 ; n682_not
g27401 not n943 ; n943_not
g27402 not n844 ; n844_not
g27403 not n754 ; n754_not
g27404 not n781 ; n781_not
g27405 not n862 ; n862_not
g27406 not n772 ; n772_not
g27407 not n961 ; n961_not
g27408 not n952 ; n952_not
g27409 not n925 ; n925_not
g27410 not n736 ; n736_not
g27411 not n727 ; n727_not
g27412 not n808 ; n808_not
g27413 not n907 ; n907_not
g27414 not n817 ; n817_not
g27415 not n763 ; n763_not
g27416 not n691 ; n691_not
g27417 not n709 ; n709_not
g27418 not n790 ; n790_not
g27419 not n826 ; n826_not
g27420 not n385 ; n385_not
g27421 not n916 ; n916_not
g27422 not n655 ; n655_not
g27423 not n646 ; n646_not
g27424 not n970 ; n970_not
g27425 not n439 ; n439_not
g27426 not n583 ; n583_not
g27427 not n448 ; n448_not
g27428 not n457 ; n457_not
g27429 not n466 ; n466_not
g27430 not n637 ; n637_not
g27431 not n475 ; n475_not
g27432 not n628 ; n628_not
g27433 not n619 ; n619_not
g27434 not n493 ; n493_not
g27435 not n529 ; n529_not
g27436 not n592 ; n592_not
g27437 not n547 ; n547_not
g27438 not n556 ; n556_not
g27439 not n565 ; n565_not
g27440 not n574 ; n574_not
g27441 not n673 ; n673_not
g27442 not n367 ; n367_not
g27443 not n358 ; n358_not
g27444 not n295 ; n295_not
g27445 not n376 ; n376_not
g27446 not n286 ; n286_not
g27447 not n664 ; n664_not
g27448 not n277 ; n277_not
g27449 not n349 ; n349_not
g27450 not n259 ; n259_not
g27451 not n890 ; n890_not
g27452 not n863 ; n863_not
g27453 not n539 ; n539_not
g27454 not n944 ; n944_not
g27455 not n908 ; n908_not
g27456 not n791 ; n791_not
g27457 not n782 ; n782_not
g27458 not n548 ; n548_not
g27459 not n773 ; n773_not
g27460 not n557 ; n557_not
g27461 not n278 ; n278_not
g27462 not n566 ; n566_not
g27463 not n575 ; n575_not
g27464 not n755 ; n755_not
g27465 not n854 ; n854_not
g27466 not n845 ; n845_not
g27467 not n926 ; n926_not
g27468 not n395 ; n395_not
g27469 not n836 ; n836_not
g27470 not n296 ; n296_not
g27471 not n827 ; n827_not
g27472 not n377 ; n377_not
g27473 not n449 ; n449_not
g27474 not n368 ; n368_not
g27475 not n458 ; n458_not
g27476 not n872 ; n872_not
g27477 not n467 ; n467_not
g27478 not n359 ; n359_not
g27479 not n881 ; n881_not
g27480 not n485 ; n485_not
g27481 not n809 ; n809_not
g27482 not n917 ; n917_not
g27483 not n764 ; n764_not
g27484 not n737 ; n737_not
g27485 not n593 ; n593_not
g27486 not n647 ; n647_not
g27487 not n728 ; n728_not
g27488 not n971 ; n971_not
g27489 not n638 ; n638_not
g27490 not n629 ; n629_not
g27491 not n719 ; n719_not
g27492 not n656 ; n656_not
g27493 not n674 ; n674_not
g27494 not n692 ; n692_not
g27495 not n962 ; n962_not
g27496 not n746 ; n746_not
g27497 not n584 ; n584_not
g27498 not n980 ; n980_not
g27499 not n819 ; n819_not
g27500 not n666 ; n666_not
g27501 not n369 ; n369_not
g27502 not n864 ; n864_not
g27503 not n486 ; n486_not
g27504 not n873 ; n873_not
g27505 not n729 ; n729_not
g27506 not n972 ; n972_not
g27507 not n918 ; n918_not
g27508 not n990 ; n990_not
g27509 not n549 ; n549_not
g27510 not n396 ; n396_not
g27511 not n657 ; n657_not
g27512 not n837 ; n837_not
g27513 not n846 ; n846_not
g27514 not n648 ; n648_not
g27515 not n828 ; n828_not
g27516 not n855 ; n855_not
g27517 not n927 ; n927_not
g27518 not n567 ; n567_not
g27519 not n954 ; n954_not
g27520 not n468 ; n468_not
g27521 not n378 ; n378_not
g27522 not n747 ; n747_not
g27523 not n792 ; n792_not
g27524 not n891 ; n891_not
g27525 not n279 ; n279_not
g27526 not n594 ; n594_not
g27527 not n765 ; n765_not
g27528 not n945 ; n945_not
g27529 not n783 ; n783_not
g27530 not n909 ; n909_not
g27531 not n459 ; n459_not
g27532 not n297 ; n297_not
g27533 not n774 ; n774_not
g27534 not n693 ; n693_not
g27535 not n936 ; n936_not
g27536 not n738 ; n738_not
g27537 not n882 ; n882_not
g27538 not n576 ; n576_not
g27539 not n675 ; n675_not
g27540 not n963 ; n963_not
g27541 not n865 ; n865_not
g27542 not n388 ; n388_not
g27543 not n667 ; n667_not
g27544 not n694 ; n694_not
g27545 not n658 ; n658_not
g27546 not n676 ; n676_not
g27547 not n685 ; n685_not
g27548 not n919 ; n919_not
g27549 not n847 ; n847_not
g27550 not n379 ; n379_not
g27551 not n964 ; n964_not
g27552 not n856 ; n856_not
g27553 not n883 ; n883_not
g27554 not n298 ; n298_not
g27555 not n874 ; n874_not
g27556 not n748 ; n748_not
g27557 not n928 ; n928_not
g27558 not n937 ; n937_not
g27559 not n496 ; n496_not
g27560 not n649 ; n649_not
g27561 not n487 ; n487_not
g27562 not n793 ; n793_not
g27563 not n478 ; n478_not
g27564 not n595 ; n595_not
g27565 not n739 ; n739_not
g27566 not n973 ; n973_not
g27567 not n469 ; n469_not
g27568 not n568 ; n568_not
g27569 not n397 ; n397_not
g27570 not n775 ; n775_not
g27571 not n838 ; n838_not
g27572 not n829 ; n829_not
g27573 not n586 ; n586_not
g27574 not n955 ; n955_not
g27575 not n938 ; n938_not
g27576 not n884 ; n884_not
g27577 not n587 ; n587_not
g27578 not n794 ; n794_not
g27579 not n983 ; n983_not
g27580 not n965 ; n965_not
g27581 not n848 ; n848_not
g27582 not n596 ; n596_not
g27583 not n299 ; n299_not
g27584 not n947 ; n947_not
g27585 not n776 ; n776_not
g27586 not n974 ; n974_not
g27587 not n686 ; n686_not
g27588 not n839 ; n839_not
g27589 not n758 ; n758_not
g27590 not n389 ; n389_not
g27591 not n398 ; n398_not
g27592 not n929 ; n929_not
g27593 not n659 ; n659_not
g27594 not n569 ; n569_not
g27595 not n857 ; n857_not
g27596 not n677 ; n677_not
g27597 not n956 ; n956_not
g27598 not n992 ; n992_not
g27599 not n668 ; n668_not
g27600 not n479 ; n479_not
g27601 not n497 ; n497_not
g27602 not n488 ; n488_not
g27603 not n875 ; n875_not
g27604 not n749 ; n749_not
g27605 not n866 ; n866_not
g27606 not n984 ; n984_not
g27607 not n993 ; n993_not
g27608 not n957 ; n957_not
g27609 not n975 ; n975_not
g27610 not n948 ; n948_not
g27611 not n966 ; n966_not
g27612 not n939 ; n939_not
g27613 not n498 ; n498_not
g27614 not n759 ; n759_not
g27615 not n849 ; n849_not
g27616 not n696 ; n696_not
g27617 not n858 ; n858_not
g27618 not n768 ; n768_not
g27619 not n867 ; n867_not
g27620 not n876 ; n876_not
g27621 not n777 ; n777_not
g27622 not n795 ; n795_not
g27623 not n687 ; n687_not
g27624 not n678 ; n678_not
g27625 not n885 ; n885_not
g27626 not n669 ; n669_not
g27627 not n579 ; n579_not
g27628 not n489 ; n489_not
g27629 not n894 ; n894_not
g27630 not n597 ; n597_not
g27631 not n588 ; n588_not
g27632 not n399 ; n399_not
g27633 not n786 ; n786_not
g27634 not n787 ; n787_not
g27635 not n967 ; n967_not
g27636 not n769 ; n769_not
g27637 not n778 ; n778_not
g27638 not n949 ; n949_not
g27639 not n679 ; n679_not
g27640 not n697 ; n697_not
g27641 not n958 ; n958_not
g27642 not n499 ; n499_not
g27643 not n976 ; n976_not
g27644 not n985 ; n985_not
g27645 not n688 ; n688_not
g27646 not n598 ; n598_not
g27647 not n589 ; n589_not
g27648 not n877 ; n877_not
g27649 not n868 ; n868_not
g27650 not n895 ; n895_not
g27651 not n796 ; n796_not
g27652 not n859 ; n859_not
g27653 not n886 ; n886_not
g27654 not n994 ; n994_not
g27655 not n878 ; n878_not
g27656 not n689 ; n689_not
g27657 not n887 ; n887_not
g27658 not n968 ; n968_not
g27659 not n896 ; n896_not
g27660 not n995 ; n995_not
g27661 not n788 ; n788_not
g27662 not n986 ; n986_not
g27663 not n779 ; n779_not
g27664 not n797 ; n797_not
g27665 not n977 ; n977_not
g27666 not n869 ; n869_not
g27667 not n959 ; n959_not
g27668 not n698 ; n698_not
g27669 not n699 ; n699_not
g27670 not n987 ; n987_not
g27671 not n996 ; n996_not
g27672 not n789 ; n789_not
g27673 not n978 ; n978_not
g27674 not n879 ; n879_not
g27675 not n897 ; n897_not
g27676 not n888 ; n888_not
g27677 not n988 ; n988_not
g27678 not n979 ; n979_not
g27679 not n997 ; n997_not
g27680 not n799 ; n799_not
g27681 not n898 ; n898_not
g27682 not n889 ; n889_not
g27683 not n998 ; n998_not
g27684 not n899 ; n899_not
g27685 not n989 ; n989_not
g27686 not n999 ; n999_not
g27687 not n1010 ; n1010_not
g27688 not n1100 ; n1100_not
g27689 not n2000 ; n2000_not
g27690 not n1101 ; n1101_not
g27691 not n1110 ; n1110_not
g27692 not n3000 ; n3000_not
g27693 not n2001 ; n2001_not
g27694 not n1002 ; n1002_not
g27695 not n1011 ; n1011_not
g27696 not n2010 ; n2010_not
g27697 not n2100 ; n2100_not
g27698 not n2101 ; n2101_not
g27699 not n2020 ; n2020_not
g27700 not n1021 ; n1021_not
g27701 not n2110 ; n2110_not
g27702 not n2011 ; n2011_not
g27703 not n2002 ; n2002_not
g27704 not n1210 ; n1210_not
g27705 not n1030 ; n1030_not
g27706 not n1120 ; n1120_not
g27707 not n3010 ; n3010_not
g27708 not n1300 ; n1300_not
g27709 not n3100 ; n3100_not
g27710 not n4000 ; n4000_not
g27711 not n1201 ; n1201_not
g27712 not n3001 ; n3001_not
g27713 not n2200 ; n2200_not
g27714 not n1111 ; n1111_not
g27715 not n1102 ; n1102_not
g27716 not n1012 ; n1012_not
g27717 not n1003 ; n1003_not
g27718 not n3110 ; n3110_not
g27719 not n3011 ; n3011_not
g27720 not n1103 ; n1103_not
g27721 not n1040 ; n1040_not
g27722 not n1301 ; n1301_not
g27723 not n4010 ; n4010_not
g27724 not n1310 ; n1310_not
g27725 not n4001 ; n4001_not
g27726 not n1004 ; n1004_not
g27727 not n2012 ; n2012_not
g27728 not n3101 ; n3101_not
g27729 not n2210 ; n2210_not
g27730 not n1202 ; n1202_not
g27731 not n1211 ; n1211_not
g27732 not n1400 ; n1400_not
g27733 not n4100 ; n4100_not
g27734 not n2021 ; n2021_not
g27735 not n2102 ; n2102_not
g27736 not n2111 ; n2111_not
g27737 not n1220 ; n1220_not
g27738 not n1013 ; n1013_not
g27739 not n2003 ; n2003_not
g27740 not n2120 ; n2120_not
g27741 not n1121 ; n1121_not
g27742 not n5000 ; n5000_not
g27743 not n1022 ; n1022_not
g27744 not n1031 ; n1031_not
g27745 not n3200 ; n3200_not
g27746 not n2030 ; n2030_not
g27747 not n1112 ; n1112_not
g27748 not n2300 ; n2300_not
g27749 not n1130 ; n1130_not
g27750 not n1221 ; n1221_not
g27751 not n1212 ; n1212_not
g27752 not n1203 ; n1203_not
g27753 not n2301 ; n2301_not
g27754 not n2310 ; n2310_not
g27755 not n5100 ; n5100_not
g27756 not n1140 ; n1140_not
g27757 not n1032 ; n1032_not
g27758 not n1122 ; n1122_not
g27759 not n2400 ; n2400_not
g27760 not n1113 ; n1113_not
g27761 not n5010 ; n5010_not
g27762 not n3300 ; n3300_not
g27763 not n3210 ; n3210_not
g27764 not n3003 ; n3003_not
g27765 not n3120 ; n3120_not
g27766 not n2013 ; n2013_not
g27767 not n2022 ; n2022_not
g27768 not n3111 ; n3111_not
g27769 not n2112 ; n2112_not
g27770 not n2121 ; n2121_not
g27771 not n2130 ; n2130_not
g27772 not n2040 ; n2040_not
g27773 not n3012 ; n3012_not
g27774 not n3102 ; n3102_not
g27775 not n3030 ; n3030_not
g27776 not n4011 ; n4011_not
g27777 not n4200 ; n4200_not
g27778 not n5001 ; n5001_not
g27779 not n1311 ; n1311_not
g27780 not n1320 ; n1320_not
g27781 not n4110 ; n4110_not
g27782 not n4101 ; n4101_not
g27783 not n1401 ; n1401_not
g27784 not n1410 ; n1410_not
g27785 not n2103 ; n2103_not
g27786 not n4020 ; n4020_not
g27787 not n4002 ; n4002_not
g27788 not n1500 ; n1500_not
g27789 not n2211 ; n2211_not
g27790 not n2220 ; n2220_not
g27791 not n1014 ; n1014_not
g27792 not n1041 ; n1041_not
g27793 not n1050 ; n1050_not
g27794 not n1023 ; n1023_not
g27795 not n1104 ; n1104_not
g27796 not n1005 ; n1005_not
g27797 not n4120 ; n4120_not
g27798 not n4201 ; n4201_not
g27799 not n3130 ; n3130_not
g27800 not n3112 ; n3112_not
g27801 not n1303 ; n1303_not
g27802 not n2113 ; n2113_not
g27803 not n3031 ; n3031_not
g27804 not n3022 ; n3022_not
g27805 not n1024 ; n1024_not
g27806 not n1312 ; n1312_not
g27807 not n5200 ; n5200_not
g27808 not n1321 ; n1321_not
g27809 not n1006 ; n1006_not
g27810 not n3121 ; n3121_not
g27811 not n1330 ; n1330_not
g27812 not n2500 ; n2500_not
g27813 not n1150 ; n1150_not
g27814 not n1204 ; n1204_not
g27815 not n3400 ; n3400_not
g27816 not n1213 ; n1213_not
g27817 not n2104 ; n2104_not
g27818 not n2041 ; n2041_not
g27819 not n1231 ; n1231_not
g27820 not n1240 ; n1240_not
g27821 not n1015 ; n1015_not
g27822 not n2203 ; n2203_not
g27823 not n2023 ; n2023_not
g27824 not n4210 ; n4210_not
g27825 not n3202 ; n3202_not
g27826 not n1600 ; n1600_not
g27827 not n4030 ; n4030_not
g27828 not n5020 ; n5020_not
g27829 not n4021 ; n4021_not
g27830 not n2140 ; n2140_not
g27831 not n4012 ; n4012_not
g27832 not n5110 ; n5110_not
g27833 not n1033 ; n1033_not
g27834 not n3211 ; n3211_not
g27835 not n6010 ; n6010_not
g27836 not n1501 ; n1501_not
g27837 not n1510 ; n1510_not
g27838 not n4003 ; n4003_not
g27839 not n3220 ; n3220_not
g27840 not n3040 ; n3040_not
g27841 not n6001 ; n6001_not
g27842 not n7000 ; n7000_not
g27843 not n6100 ; n6100_not
g27844 not n4111 ; n4111_not
g27845 not n2302 ; n2302_not
g27846 not n4102 ; n4102_not
g27847 not n1402 ; n1402_not
g27848 not n1411 ; n1411_not
g27849 not n3301 ; n3301_not
g27850 not n2122 ; n2122_not
g27851 not n5101 ; n5101_not
g27852 not n1420 ; n1420_not
g27853 not n2311 ; n2311_not
g27854 not n1042 ; n1042_not
g27855 not n2410 ; n2410_not
g27856 not n2131 ; n2131_not
g27857 not n2401 ; n2401_not
g27858 not n3013 ; n3013_not
g27859 not n1141 ; n1141_not
g27860 not n3004 ; n3004_not
g27861 not n1132 ; n1132_not
g27862 not n2014 ; n2014_not
g27863 not n3103 ; n3103_not
g27864 not n2221 ; n2221_not
g27865 not n2212 ; n2212_not
g27866 not n1114 ; n1114_not
g27867 not n1105 ; n1105_not
g27868 not n1051 ; n1051_not
g27869 not n4300 ; n4300_not
g27870 not n5011 ; n5011_not
g27871 not n5002 ; n5002_not
g27872 not n2230 ; n2230_not
g27873 not n3104 ; n3104_not
g27874 not n3131 ; n3131_not
g27875 not n2141 ; n2141_not
g27876 not n3140 ; n3140_not
g27877 not n4121 ; n4121_not
g27878 not n3005 ; n3005_not
g27879 not n4112 ; n4112_not
g27880 not n6101 ; n6101_not
g27881 not n1322 ; n1322_not
g27882 not n4301 ; n4301_not
g27883 not n2303 ; n2303_not
g27884 not n2231 ; n2231_not
g27885 not n4103 ; n4103_not
g27886 not n1061 ; n1061_not
g27887 not n1070 ; n1070_not
g27888 not n1403 ; n1403_not
g27889 not n3302 ; n3302_not
g27890 not n4130 ; n4130_not
g27891 not n1412 ; n1412_not
g27892 not n5210 ; n5210_not
g27893 not n2006 ; n2006_not
g27894 not n1025 ; n1025_not
g27895 not n5201 ; n5201_not
g27896 not n6200 ; n6200_not
g27897 not n1313 ; n1313_not
g27898 not n1160 ; n1160_not
g27899 not n3122 ; n3122_not
g27900 not n4310 ; n4310_not
g27901 not n3023 ; n3023_not
g27902 not n1331 ; n1331_not
g27903 not n3113 ; n3113_not
g27904 not n1151 ; n1151_not
g27905 not n4040 ; n4040_not
g27906 not n2051 ; n2051_not
g27907 not n1340 ; n1340_not
g27908 not n3032 ; n3032_not
g27909 not n5012 ; n5012_not
g27910 not n4400 ; n4400_not
g27911 not n2132 ; n2132_not
g27912 not n3320 ; n3320_not
g27913 not n2222 ; n2222_not
g27914 not n6011 ; n6011_not
g27915 not n1115 ; n1115_not
g27916 not n1052 ; n1052_not
g27917 not n1502 ; n1502_not
g27918 not n3212 ; n3212_not
g27919 not n4004 ; n4004_not
g27920 not n1511 ; n1511_not
g27921 not n6110 ; n6110_not
g27922 not n5111 ; n5111_not
g27923 not n3221 ; n3221_not
g27924 not n1520 ; n1520_not
g27925 not n1421 ; n1421_not
g27926 not n6002 ; n6002_not
g27927 not n5120 ; n5120_not
g27928 not n1106 ; n1106_not
g27929 not n7010 ; n7010_not
g27930 not n3041 ; n3041_not
g27931 not n2150 ; n2150_not
g27932 not n7100 ; n7100_not
g27933 not n5003 ; n5003_not
g27934 not n2420 ; n2420_not
g27935 not n2123 ; n2123_not
g27936 not n1430 ; n1430_not
g27937 not n1133 ; n1133_not
g27938 not n2312 ; n2312_not
g27939 not n1043 ; n1043_not
g27940 not n5102 ; n5102_not
g27941 not n2411 ; n2411_not
g27942 not n5021 ; n5021_not
g27943 not n2321 ; n2321_not
g27944 not n3014 ; n3014_not
g27945 not n1601 ; n1601_not
g27946 not n2402 ; n2402_not
g27947 not n6020 ; n6020_not
g27948 not n2330 ; n2330_not
g27949 not n4022 ; n4022_not
g27950 not n3203 ; n3203_not
g27951 not n2033 ; n2033_not
g27952 not n1007 ; n1007_not
g27953 not n8000 ; n8000_not
g27954 not n3500 ; n3500_not
g27955 not n3410 ; n3410_not
g27956 not n2015 ; n2015_not
g27957 not n2204 ; n2204_not
g27958 not n4220 ; n4220_not
g27959 not n1250 ; n1250_not
g27960 not n3401 ; n3401_not
g27961 not n2240 ; n2240_not
g27962 not n1205 ; n1205_not
g27963 not n1223 ; n1223_not
g27964 not n2024 ; n2024_not
g27965 not n2105 ; n2105_not
g27966 not n1016 ; n1016_not
g27967 not n2501 ; n2501_not
g27968 not n2042 ; n2042_not
g27969 not n4202 ; n4202_not
g27970 not n5300 ; n5300_not
g27971 not n1241 ; n1241_not
g27972 not n2213 ; n2213_not
g27973 not n4211 ; n4211_not
g27974 not n1232 ; n1232_not
g27975 not n2060 ; n2060_not
g27976 not n2403 ; n2403_not
g27977 not n1125 ; n1125_not
g27978 not n1620 ; n1620_not
g27979 not n5211 ; n5211_not
g27980 not n4320 ; n4320_not
g27981 not n7200 ; n7200_not
g27982 not n2322 ; n2322_not
g27983 not n1602 ; n1602_not
g27984 not n4050 ; n4050_not
g27985 not n5301 ; n5301_not
g27986 not n3240 ; n3240_not
g27987 not n2223 ; n2223_not
g27988 not n5022 ; n5022_not
g27989 not n1413 ; n1413_not
g27990 not n3105 ; n3105_not
g27991 not n1404 ; n1404_not
g27992 not n3042 ; n3042_not
g27993 not n1107 ; n1107_not
g27994 not n8100 ; n8100_not
g27995 not n3501 ; n3501_not
g27996 not n5013 ; n5013_not
g27997 not n1233 ; n1233_not
g27998 not n3150 ; n3150_not
g27999 not n1134 ; n1134_not
g28000 not n1422 ; n1422_not
g28001 not n2124 ; n2124_not
g28002 not n4230 ; n4230_not
g28003 not n1431 ; n1431_not
g28004 not n2106 ; n2106_not
g28005 not n2313 ; n2313_not
g28006 not n2412 ; n2412_not
g28007 not n4122 ; n4122_not
g28008 not n1440 ; n1440_not
g28009 not n2610 ; n2610_not
g28010 not n1305 ; n1305_not
g28011 not n6021 ; n6021_not
g28012 not n2142 ; n2142_not
g28013 not n6111 ; n6111_not
g28014 not n5031 ; n5031_not
g28015 not n1161 ; n1161_not
g28016 not n1521 ; n1521_not
g28017 not n5130 ; n5130_not
g28018 not n6003 ; n6003_not
g28019 not n2214 ; n2214_not
g28020 not n2340 ; n2340_not
g28021 not n3222 ; n3222_not
g28022 not n2052 ; n2052_not
g28023 not n5112 ; n5112_not
g28024 not n7020 ; n7020_not
g28025 not n5121 ; n5121_not
g28026 not n7011 ; n7011_not
g28027 not n3510 ; n3510_not
g28028 not n7101 ; n7101_not
g28029 not n3060 ; n3060_not
g28030 not n2151 ; n2151_not
g28031 not n2133 ; n2133_not
g28032 not n2502 ; n2502_not
g28033 not n2241 ; n2241_not
g28034 not n2205 ; n2205_not
g28035 not n3051 ; n3051_not
g28036 not n4023 ; n4023_not
g28037 not n2511 ; n2511_not
g28038 not n1215 ; n1215_not
g28039 not n4410 ; n4410_not
g28040 not n3204 ; n3204_not
g28041 not n2160 ; n2160_not
g28042 not n4014 ; n4014_not
g28043 not n4104 ; n4104_not
g28044 not n4221 ; n4221_not
g28045 not n1080 ; n1080_not
g28046 not n2601 ; n2601_not
g28047 not n1035 ; n1035_not
g28048 not n1053 ; n1053_not
g28049 not n2250 ; n2250_not
g28050 not n1116 ; n1116_not
g28051 not n1503 ; n1503_not
g28052 not n1512 ; n1512_not
g28053 not n1017 ; n1017_not
g28054 not n2025 ; n2025_not
g28055 not n1323 ; n1323_not
g28056 not n3123 ; n3123_not
g28057 not n4212 ; n4212_not
g28058 not n1332 ; n1332_not
g28059 not n6201 ; n6201_not
g28060 not n6210 ; n6210_not
g28061 not n1341 ; n1341_not
g28062 not n4140 ; n4140_not
g28063 not n3321 ; n3321_not
g28064 not n1350 ; n1350_not
g28065 not n5040 ; n5040_not
g28066 not n2700 ; n2700_not
g28067 not n4131 ; n4131_not
g28068 not n5310 ; n5310_not
g28069 not n4041 ; n4041_not
g28070 not n1152 ; n1152_not
g28071 not n5004 ; n5004_not
g28072 not n7110 ; n7110_not
g28073 not n2520 ; n2520_not
g28074 not n2016 ; n2016_not
g28075 not n3213 ; n3213_not
g28076 not n5220 ; n5220_not
g28077 not n3114 ; n3114_not
g28078 not n1071 ; n1071_not
g28079 not n3411 ; n3411_not
g28080 not n2070 ; n2070_not
g28081 not n4203 ; n4203_not
g28082 not n3600 ; n3600_not
g28083 not n3024 ; n3024_not
g28084 not n2007 ; n2007_not
g28085 not n1314 ; n1314_not
g28086 not n1170 ; n1170_not
g28087 not n3015 ; n3015_not
g28088 not n4302 ; n4302_not
g28089 not n5202 ; n5202_not
g28090 not n3420 ; n3420_not
g28091 not n2421 ; n2421_not
g28092 not n3006 ; n3006_not
g28093 not n2430 ; n2430_not
g28094 not n6120 ; n6120_not
g28095 not n3141 ; n3141_not
g28096 not n1251 ; n1251_not
g28097 not n6030 ; n6030_not
g28098 not n2115 ; n2115_not
g28099 not n1062 ; n1062_not
g28100 not n3303 ; n3303_not
g28101 not n2034 ; n2034_not
g28102 not n2232 ; n2232_not
g28103 not n1242 ; n1242_not
g28104 not n2304 ; n2304_not
g28105 not n2061 ; n2061_not
g28106 not n8010 ; n8010_not
g28107 not n4500 ; n4500_not
g28108 not n1710 ; n1710_not
g28109 not n3312 ; n3312_not
g28110 not n5113 ; n5113_not
g28111 not n3520 ; n3520_not
g28112 not n2323 ; n2323_not
g28113 not n3250 ; n3250_not
g28114 not n5302 ; n5302_not
g28115 not n1603 ; n1603_not
g28116 not n1801 ; n1801_not
g28117 not n3313 ; n3313_not
g28118 not n5320 ; n5320_not
g28119 not n6400 ; n6400_not
g28120 not n1630 ; n1630_not
g28121 not n7102 ; n7102_not
g28122 not n2233 ; n2233_not
g28123 not n6004 ; n6004_not
g28124 not n3340 ; n3340_not
g28125 not n5014 ; n5014_not
g28126 not n2341 ; n2341_not
g28127 not n3412 ; n3412_not
g28128 not n2242 ; n2242_not
g28129 not n1900 ; n1900_not
g28130 not n7300 ; n7300_not
g28131 not n6112 ; n6112_not
g28132 not n1612 ; n1612_not
g28133 not n8101 ; n8101_not
g28134 not n3601 ; n3601_not
g28135 not n3430 ; n3430_not
g28136 not n3700 ; n3700_not
g28137 not n2224 ; n2224_not
g28138 not n3610 ; n3610_not
g28139 not n1036 ; n1036_not
g28140 not n2152 ; n2152_not
g28141 not n5041 ; n5041_not
g28142 not n2305 ; n2305_not
g28143 not n3421 ; n3421_not
g28144 not n5023 ; n5023_not
g28145 not n4600 ; n4600_not
g28146 not n3241 ; n3241_not
g28147 not n2143 ; n2143_not
g28148 not n6310 ; n6310_not
g28149 not n2206 ; n2206_not
g28150 not n1711 ; n1711_not
g28151 not n2260 ; n2260_not
g28152 not n1810 ; n1810_not
g28153 not n3322 ; n3322_not
g28154 not n6040 ; n6040_not
g28155 not n3043 ; n3043_not
g28156 not n2161 ; n2161_not
g28157 not n1702 ; n1702_not
g28158 not n3502 ; n3502_not
g28159 not n1522 ; n1522_not
g28160 not n3331 ; n3331_not
g28161 not n1540 ; n1540_not
g28162 not n2251 ; n2251_not
g28163 not n5032 ; n5032_not
g28164 not n1720 ; n1720_not
g28165 not n5050 ; n5050_not
g28166 not n8110 ; n8110_not
g28167 not n6022 ; n6022_not
g28168 not n8011 ; n8011_not
g28169 not n3304 ; n3304_not
g28170 not n3214 ; n3214_not
g28171 not n8020 ; n8020_not
g28172 not n8200 ; n8200_not
g28173 not n1621 ; n1621_not
g28174 not n2170 ; n2170_not
g28175 not n3025 ; n3025_not
g28176 not n4312 ; n4312_not
g28177 not n2008 ; n2008_not
g28178 not n1306 ; n1306_not
g28179 not n6121 ; n6121_not
g28180 not n1072 ; n1072_not
g28181 not n3115 ; n3115_not
g28182 not n4510 ; n4510_not
g28183 not n1018 ; n1018_not
g28184 not n5221 ; n5221_not
g28185 not n4204 ; n4204_not
g28186 not n2017 ; n2017_not
g28187 not n4213 ; n4213_not
g28188 not n4501 ; n4501_not
g28189 not n1270 ; n1270_not
g28190 not n4222 ; n4222_not
g28191 not n2026 ; n2026_not
g28192 not n5311 ; n5311_not
g28193 not n2620 ; n2620_not
g28194 not n5230 ; n5230_not
g28195 not n7111 ; n7111_not
g28196 not n1009 ; n1009_not
g28197 not n1324 ; n1324_not
g28198 not n3142 ; n3142_not
g28199 not n2431 ; n2431_not
g28200 not n3133 ; n3133_not
g28201 not n4123 ; n4123_not
g28202 not n2701 ; n2701_not
g28203 not n2116 ; n2116_not
g28204 not n1360 ; n1360_not
g28205 not n4132 ; n4132_not
g28206 not n6220 ; n6220_not
g28207 not n1351 ; n1351_not
g28208 not n4141 ; n4141_not
g28209 not n3124 ; n3124_not
g28210 not n5410 ; n5410_not
g28211 not n1342 ; n1342_not
g28212 not n1225 ; n1225_not
g28213 not n1243 ; n1243_not
g28214 not n2440 ; n2440_not
g28215 not n1333 ; n1333_not
g28216 not n9100 ; n9100_not
g28217 not n5203 ; n5203_not
g28218 not n1315 ; n1315_not
g28219 not n2512 ; n2512_not
g28220 not n2062 ; n2062_not
g28221 not n1090 ; n1090_not
g28222 not n1171 ; n1171_not
g28223 not n7120 ; n7120_not
g28224 not n1162 ; n1162_not
g28225 not n2521 ; n2521_not
g28226 not n4303 ; n4303_not
g28227 not n1153 ; n1153_not
g28228 not n4240 ; n4240_not
g28229 not n2530 ; n2530_not
g28230 not n2071 ; n2071_not
g28231 not n1144 ; n1144_not
g28232 not n7012 ; n7012_not
g28233 not n4330 ; n4330_not
g28234 not n1135 ; n1135_not
g28235 not n1126 ; n1126_not
g28236 not n2080 ; n2080_not
g28237 not n4321 ; n4321_not
g28238 not n1108 ; n1108_not
g28239 not n1252 ; n1252_not
g28240 not n4231 ; n4231_not
g28241 not n2035 ; n2035_not
g28242 not n1234 ; n1234_not
g28243 not n2611 ; n2611_not
g28244 not n2107 ; n2107_not
g28245 not n2602 ; n2602_not
g28246 not n6031 ; n6031_not
g28247 not n2503 ; n2503_not
g28248 not n2044 ; n2044_not
g28249 not n1207 ; n1207_not
g28250 not n1081 ; n1081_not
g28251 not n2053 ; n2053_not
g28252 not n6202 ; n6202_not
g28253 not n6130 ; n6130_not
g28254 not n3106 ; n3106_not
g28255 not n1180 ; n1180_not
g28256 not n4024 ; n4024_not
g28257 not n2134 ; n2134_not
g28258 not n4033 ; n4033_not
g28259 not n1450 ; n1450_not
g28260 not n7210 ; n7210_not
g28261 not n3070 ; n3070_not
g28262 not n4042 ; n4042_not
g28263 not n2404 ; n2404_not
g28264 not n4051 ; n4051_not
g28265 not n3016 ; n3016_not
g28266 not n4060 ; n4060_not
g28267 not n3151 ; n3151_not
g28268 not n2350 ; n2350_not
g28269 not n5212 ; n5212_not
g28270 not n1441 ; n1441_not
g28271 not n7003 ; n7003_not
g28272 not n3061 ; n3061_not
g28273 not n3232 ; n3232_not
g28274 not n3223 ; n3223_not
g28275 not n5122 ; n5122_not
g28276 not n1531 ; n1531_not
g28277 not n2800 ; n2800_not
g28278 not n9010 ; n9010_not
g28279 not n7021 ; n7021_not
g28280 not n1504 ; n1504_not
g28281 not n1513 ; n1513_not
g28282 not n5131 ; n5131_not
g28283 not n5140 ; n5140_not
g28284 not n3205 ; n3205_not
g28285 not n4015 ; n4015_not
g28286 not n1405 ; n1405_not
g28287 not n2422 ; n2422_not
g28288 not n1414 ; n1414_not
g28289 not n1054 ; n1054_not
g28290 not n1063 ; n1063_not
g28291 not n4105 ; n4105_not
g28292 not n7030 ; n7030_not
g28293 not n2710 ; n2710_not
g28294 not n2125 ; n2125_not
g28295 not n1432 ; n1432_not
g28296 not n1423 ; n1423_not
g28297 not n7201 ; n7201_not
g28298 not n3160 ; n3160_not
g28299 not n2063 ; n2063_not
g28300 not n2027 ; n2027_not
g28301 not n2144 ; n2144_not
g28302 not n2081 ; n2081_not
g28303 not n3314 ; n3314_not
g28304 not n3251 ; n3251_not
g28305 not n1802 ; n1802_not
g28306 not n5420 ; n5420_not
g28307 not n3107 ; n3107_not
g28308 not n3053 ; n3053_not
g28309 not n2054 ; n2054_not
g28310 not n3215 ; n3215_not
g28311 not n7022 ; n7022_not
g28312 not n2090 ; n2090_not
g28313 not n3125 ; n3125_not
g28314 not n3404 ; n3404_not
g28315 not n6113 ; n6113_not
g28316 not n6410 ; n6410_not
g28317 not n1910 ; n1910_not
g28318 not n3233 ; n3233_not
g28319 not n3305 ; n3305_not
g28320 not n2153 ; n2153_not
g28321 not n3143 ; n3143_not
g28322 not n3080 ; n3080_not
g28323 not n9200 ; n9200_not
g28324 not n3224 ; n3224_not
g28325 not n5015 ; n5015_not
g28326 not n1901 ; n1901_not
g28327 not n2117 ; n2117_not
g28328 not n3062 ; n3062_not
g28329 not n9020 ; n9020_not
g28330 not n3413 ; n3413_not
g28331 not n3134 ; n3134_not
g28332 not n3071 ; n3071_not
g28333 not n3332 ; n3332_not
g28334 not n6104 ; n6104_not
g28335 not n8102 ; n8102_not
g28336 not n3170 ; n3170_not
g28337 not n3026 ; n3026_not
g28338 not n1820 ; n1820_not
g28339 not n8120 ; n8120_not
g28340 not n3152 ; n3152_not
g28341 not n1019 ; n1019_not
g28342 not n6302 ; n6302_not
g28343 not n6131 ; n6131_not
g28344 not n3044 ; n3044_not
g28345 not n2171 ; n2171_not
g28346 not n7103 ; n7103_not
g28347 not n2126 ; n2126_not
g28348 not n3017 ; n3017_not
g28349 not n3116 ; n3116_not
g28350 not n2009 ; n2009_not
g28351 not n3350 ; n3350_not
g28352 not n3341 ; n3341_not
g28353 not n3161 ; n3161_not
g28354 not n1037 ; n1037_not
g28355 not n6122 ; n6122_not
g28356 not n5510 ; n5510_not
g28357 not n5411 ; n5411_not
g28358 not n3323 ; n3323_not
g28359 not n1811 ; n1811_not
g28360 not n3035 ; n3035_not
g28361 not n4403 ; n4403_not
g28362 not n2207 ; n2207_not
g28363 not n2045 ; n2045_not
g28364 not n5402 ; n5402_not
g28365 not n6401 ; n6401_not
g28366 not n1028 ; n1028_not
g28367 not n6032 ; n6032_not
g28368 not n6320 ; n6320_not
g28369 not n9110 ; n9110_not
g28370 not n2036 ; n2036_not
g28371 not n6311 ; n6311_not
g28372 not n2135 ; n2135_not
g28373 not n2108 ; n2108_not
g28374 not n1064 ; n1064_not
g28375 not n6221 ; n6221_not
g28376 not n2711 ; n2711_not
g28377 not n1316 ; n1316_not
g28378 not n4106 ; n4106_not
g28379 not n1406 ; n1406_not
g28380 not n1415 ; n1415_not
g28381 not n2423 ; n2423_not
g28382 not n2720 ; n2720_not
g28383 not n1424 ; n1424_not
g28384 not n2414 ; n2414_not
g28385 not n1433 ; n1433_not
g28386 not n4070 ; n4070_not
g28387 not n7202 ; n7202_not
g28388 not n1442 ; n1442_not
g28389 not n4061 ; n4061_not
g28390 not n2441 ; n2441_not
g28391 not n1334 ; n1334_not
g28392 not n1244 ; n1244_not
g28393 not n4133 ; n4133_not
g28394 not n1343 ; n1343_not
g28395 not n4142 ; n4142_not
g28396 not n1235 ; n1235_not
g28397 not n1352 ; n1352_not
g28398 not n1361 ; n1361_not
g28399 not n4052 ; n4052_not
g28400 not n4124 ; n4124_not
g28401 not n1370 ; n1370_not
g28402 not n2432 ; n2432_not
g28403 not n4115 ; n4115_not
g28404 not n4007 ; n4007_not
g28405 not n5141 ; n5141_not
g28406 not n5132 ; n5132_not
g28407 not n1505 ; n1505_not
g28408 not n1514 ; n1514_not
g28409 not n9011 ; n9011_not
g28410 not n1046 ; n1046_not
g28411 not n7220 ; n7220_not
g28412 not n1523 ; n1523_not
g28413 not n1532 ; n1532_not
g28414 not n2810 ; n2810_not
g28415 not n7013 ; n7013_not
g28416 not n1541 ; n1541_not
g28417 not n7112 ; n7112_not
g28418 not n2360 ; n2360_not
g28419 not n6230 ; n6230_not
g28420 not n1451 ; n1451_not
g28421 not n2405 ; n2405_not
g28422 not n2351 ; n2351_not
g28423 not n4043 ; n4043_not
g28424 not n7211 ; n7211_not
g28425 not n1460 ; n1460_not
g28426 not n4034 ; n4034_not
g28427 not n5330 ; n5330_not
g28428 not n9002 ; n9002_not
g28429 not n5150 ; n5150_not
g28430 not n4016 ; n4016_not
g28431 not n1181 ; n1181_not
g28432 not n2504 ; n2504_not
g28433 not n4331 ; n4331_not
g28434 not n1190 ; n1190_not
g28435 not n1172 ; n1172_not
g28436 not n4250 ; n4250_not
g28437 not n1082 ; n1082_not
g28438 not n7040 ; n7040_not
g28439 not n4241 ; n4241_not
g28440 not n2603 ; n2603_not
g28441 not n1217 ; n1217_not
g28442 not n1109 ; n1109_not
g28443 not n1118 ; n1118_not
g28444 not n2531 ; n2531_not
g28445 not n4313 ; n4313_not
g28446 not n4322 ; n4322_not
g28447 not n1127 ; n1127_not
g28448 not n5051 ; n5051_not
g28449 not n1136 ; n1136_not
g28450 not n2540 ; n2540_not
g28451 not n1145 ; n1145_not
g28452 not n1091 ; n1091_not
g28453 not n4304 ; n4304_not
g28454 not n1163 ; n1163_not
g28455 not n7121 ; n7121_not
g28456 not n2513 ; n2513_not
g28457 not n6203 ; n6203_not
g28458 not n4205 ; n4205_not
g28459 not n5222 ; n5222_not
g28460 not n4511 ; n4511_not
g28461 not n5213 ; n5213_not
g28462 not n1307 ; n1307_not
g28463 not n5321 ; n5321_not
g28464 not n7031 ; n7031_not
g28465 not n5204 ; n5204_not
g28466 not n1325 ; n1325_not
g28467 not n2315 ; n2315_not
g28468 not n4160 ; n4160_not
g28469 not n4151 ; n4151_not
g28470 not n4340 ; n4340_not
g28471 not n1226 ; n1226_not
g28472 not n5303 ; n5303_not
g28473 not n4232 ; n4232_not
g28474 not n5231 ; n5231_not
g28475 not n1253 ; n1253_not
g28476 not n1262 ; n1262_not
g28477 not n2621 ; n2621_not
g28478 not n1271 ; n1271_not
g28479 not n4214 ; n4214_not
g28480 not n2630 ; n2630_not
g28481 not n1280 ; n1280_not
g28482 not n8030 ; n8030_not
g28483 not n6050 ; n6050_not
g28484 not n3611 ; n3611_not
g28485 not n5042 ; n5042_not
g28486 not n3620 ; n3620_not
g28487 not n2270 ; n2270_not
g28488 not n6041 ; n6041_not
g28489 not n5060 ; n5060_not
g28490 not n7310 ; n7310_not
g28491 not n3602 ; n3602_not
g28492 not n3701 ; n3701_not
g28493 not n3710 ; n3710_not
g28494 not n2900 ; n2900_not
g28495 not n8300 ; n8300_not
g28496 not n1604 ; n1604_not
g28497 not n4700 ; n4700_not
g28498 not n1640 ; n1640_not
g28499 not n2306 ; n2306_not
g28500 not n3800 ; n3800_not
g28501 not n1631 ; n1631_not
g28502 not n4502 ; n4502_not
g28503 not n6023 ; n6023_not
g28504 not n3431 ; n3431_not
g28505 not n4430 ; n4430_not
g28506 not n4412 ; n4412_not
g28507 not n3440 ; n3440_not
g28508 not n3422 ; n3422_not
g28509 not n5024 ; n5024_not
g28510 not n8021 ; n8021_not
g28511 not n8012 ; n8012_not
g28512 not n3503 ; n3503_not
g28513 not n2243 ; n2243_not
g28514 not n3512 ; n3512_not
g28515 not n3521 ; n3521_not
g28516 not n5033 ; n5033_not
g28517 not n1730 ; n1730_not
g28518 not n2252 ; n2252_not
g28519 not n3530 ; n3530_not
g28520 not n2180 ; n2180_not
g28521 not n1721 ; n1721_not
g28522 not n8201 ; n8201_not
g28523 not n8003 ; n8003_not
g28524 not n1712 ; n1712_not
g28525 not n6500 ; n6500_not
g28526 not n1703 ; n1703_not
g28527 not n8210 ; n8210_not
g28528 not n4610 ; n4610_not
g28529 not n6005 ; n6005_not
g28530 not n2342 ; n2342_not
g28531 not n4601 ; n4601_not
g28532 not n5600 ; n5600_not
g28533 not n5114 ; n5114_not
g28534 not n6014 ; n6014_not
g28535 not n7301 ; n7301_not
g28536 not n2333 ; n2333_not
g28537 not n7004 ; n7004_not
g28538 not n2324 ; n2324_not
g28539 not n1613 ; n1613_not
g28540 not n5105 ; n5105_not
g28541 not n1550 ; n1550_not
g28542 not n2801 ; n2801_not
g28543 not n7400 ; n7400_not
g28544 not n3081 ; n3081_not
g28545 not n8400 ; n8400_not
g28546 not n5232 ; n5232_not
g28547 not n3063 ; n3063_not
g28548 not n5115 ; n5115_not
g28549 not n5151 ; n5151_not
g28550 not n6240 ; n6240_not
g28551 not n2532 ; n2532_not
g28552 not n5331 ; n5331_not
g28553 not n2604 ; n2604_not
g28554 not n5034 ; n5034_not
g28555 not n2820 ; n2820_not
g28556 not n2811 ; n2811_not
g28557 not n9003 ; n9003_not
g28558 not n2262 ; n2262_not
g28559 not n4431 ; n4431_not
g28560 not n5304 ; n5304_not
g28561 not n8211 ; n8211_not
g28562 not n3018 ; n3018_not
g28563 not n3090 ; n3090_not
g28564 not n3009 ; n3009_not
g28565 not n2352 ; n2352_not
g28566 not n5340 ; n5340_not
g28567 not n4422 ; n4422_not
g28568 not n3072 ; n3072_not
g28569 not n2550 ; n2550_not
g28570 not n5061 ; n5061_not
g28571 not n2217 ; n2217_not
g28572 not n2505 ; n2505_not
g28573 not n2361 ; n2361_not
g28574 not n5250 ; n5250_not
g28575 not n2514 ; n2514_not
g28576 not n2226 ; n2226_not
g28577 not n2370 ; n2370_not
g28578 not n2244 ; n2244_not
g28579 not n2802 ; n2802_not
g28580 not n2208 ; n2208_not
g28581 not n2091 ; n2091_not
g28582 not n6006 ; n6006_not
g28583 not n8031 ; n8031_not
g28584 not n8202 ; n8202_not
g28585 not n9012 ; n9012_not
g28586 not n2181 ; n2181_not
g28587 not n2325 ; n2325_not
g28588 not n2433 ; n2433_not
g28589 not n3036 ; n3036_not
g28590 not n2901 ; n2901_not
g28591 not n2910 ; n2910_not
g28592 not n9030 ; n9030_not
g28593 not n5070 ; n5070_not
g28594 not n6141 ; n6141_not
g28595 not n6123 ; n6123_not
g28596 not n5205 ; n5205_not
g28597 not n2730 ; n2730_not
g28598 not n6213 ; n6213_not
g28599 not n5106 ; n5106_not
g28600 not n2334 ; n2334_not
g28601 not n2172 ; n2172_not
g28602 not n2316 ; n2316_not
g28603 not n2415 ; n2415_not
g28604 not n6222 ; n6222_not
g28605 not n2127 ; n2127_not
g28606 not n2307 ; n2307_not
g28607 not n2424 ; n2424_not
g28608 not n4404 ; n4404_not
g28609 not n2406 ; n2406_not
g28610 not n6132 ; n6132_not
g28611 not n4413 ; n4413_not
g28612 not n8310 ; n8310_not
g28613 not n5016 ; n5016_not
g28614 not n2460 ; n2460_not
g28615 not n5025 ; n5025_not
g28616 not n2640 ; n2640_not
g28617 not n2271 ; n2271_not
g28618 not n8220 ; n8220_not
g28619 not n2190 ; n2190_not
g28620 not n3027 ; n3027_not
g28621 not n2631 ; n2631_not
g28622 not n5043 ; n5043_not
g28623 not n2154 ; n2154_not
g28624 not n2622 ; n2622_not
g28625 not n2064 ; n2064_not
g28626 not n5160 ; n5160_not
g28627 not n2109 ; n2109_not
g28628 not n2442 ; n2442_not
g28629 not n2280 ; n2280_not
g28630 not n6150 ; n6150_not
g28631 not n5052 ; n5052_not
g28632 not n5322 ; n5322_not
g28633 not n2136 ; n2136_not
g28634 not n6204 ; n6204_not
g28635 not n5214 ; n5214_not
g28636 not n3054 ; n3054_not
g28637 not n5610 ; n5610_not
g28638 not n7005 ; n7005_not
g28639 not n1551 ; n1551_not
g28640 not n7302 ; n7302_not
g28641 not n1560 ; n1560_not
g28642 not n5601 ; n5601_not
g28643 not n4602 ; n4602_not
g28644 not n7320 ; n7320_not
g28645 not n3900 ; n3900_not
g28646 not n7050 ; n7050_not
g28647 not n4350 ; n4350_not
g28648 not n4611 ; n4611_not
g28649 not n6015 ; n6015_not
g28650 not n7401 ; n7401_not
g28651 not n1605 ; n1605_not
g28652 not n1614 ; n1614_not
g28653 not n4503 ; n4503_not
g28654 not n4035 ; n4035_not
g28655 not n1470 ; n1470_not
g28656 not n4026 ; n4026_not
g28657 not n4017 ; n4017_not
g28658 not n1047 ; n1047_not
g28659 not n4008 ; n4008_not
g28660 not n7212 ; n7212_not
g28661 not n7203 ; n7203_not
g28662 not n1506 ; n1506_not
g28663 not n1515 ; n1515_not
g28664 not n1524 ; n1524_not
g28665 not n7230 ; n7230_not
g28666 not n7221 ; n7221_not
g28667 not n1533 ; n1533_not
g28668 not n7014 ; n7014_not
g28669 not n1542 ; n1542_not
g28670 not n3630 ; n3630_not
g28671 not n3612 ; n3612_not
g28672 not n6051 ; n6051_not
g28673 not n3603 ; n3603_not
g28674 not n6510 ; n6510_not
g28675 not n6501 ; n6501_not
g28676 not n1704 ; n1704_not
g28677 not n1713 ; n1713_not
g28678 not n8004 ; n8004_not
g28679 not n3540 ; n3540_not
g28680 not n6060 ; n6060_not
g28681 not n3531 ; n3531_not
g28682 not n3342 ; n3342_not
g28683 not n1731 ; n1731_not
g28684 not n3522 ; n3522_not
g28685 not n1740 ; n1740_not
g28686 not n3513 ; n3513_not
g28687 not n1623 ; n1623_not
g28688 not n1632 ; n1632_not
g28689 not n3801 ; n3801_not
g28690 not n7500 ; n7500_not
g28691 not n7410 ; n7410_not
g28692 not n1641 ; n1641_not
g28693 not n4701 ; n4701_not
g28694 not n4710 ; n4710_not
g28695 not n1650 ; n1650_not
g28696 not n3504 ; n3504_not
g28697 not n3720 ; n3720_not
g28698 not n3702 ; n3702_not
g28699 not n6033 ; n6033_not
g28700 not n6600 ; n6600_not
g28701 not n1038 ; n1038_not
g28702 not n4800 ; n4800_not
g28703 not n6042 ; n6042_not
g28704 not n7041 ; n7041_not
g28705 not n1209 ; n1209_not
g28706 not n4332 ; n4332_not
g28707 not n1137 ; n1137_not
g28708 not n1218 ; n1218_not
g28709 not n4242 ; n4242_not
g28710 not n1119 ; n1119_not
g28711 not n4341 ; n4341_not
g28712 not n1227 ; n1227_not
g28713 not n4233 ; n4233_not
g28714 not n1236 ; n1236_not
g28715 not n1245 ; n1245_not
g28716 not n1254 ; n1254_not
g28717 not n1263 ; n1263_not
g28718 not n4224 ; n4224_not
g28719 not n4314 ; n4314_not
g28720 not n1128 ; n1128_not
g28721 not n4251 ; n4251_not
g28722 not n1146 ; n1146_not
g28723 not n4305 ; n4305_not
g28724 not n1164 ; n1164_not
g28725 not n7113 ; n7113_not
g28726 not n1173 ; n1173_not
g28727 not n7122 ; n7122_not
g28728 not n5511 ; n5511_not
g28729 not n1182 ; n1182_not
g28730 not n7140 ; n7140_not
g28731 not n4260 ; n4260_not
g28732 not n1191 ; n1191_not
g28733 not n5700 ; n5700_not
g28734 not n4134 ; n4134_not
g28735 not n4125 ; n4125_not
g28736 not n1371 ; n1371_not
g28737 not n4116 ; n4116_not
g28738 not n4107 ; n4107_not
g28739 not n4053 ; n4053_not
g28740 not n1407 ; n1407_not
g28741 not n1416 ; n1416_not
g28742 not n4530 ; n4530_not
g28743 not n4071 ; n4071_not
g28744 not n1425 ; n1425_not
g28745 not n4080 ; n4080_not
g28746 not n1434 ; n1434_not
g28747 not n1443 ; n1443_not
g28748 not n4062 ; n4062_not
g28749 not n1362 ; n1362_not
g28750 not n7023 ; n7023_not
g28751 not n4044 ; n4044_not
g28752 not n4206 ; n4206_not
g28753 not n1290 ; n1290_not
g28754 not n7032 ; n7032_not
g28755 not n4512 ; n4512_not
g28756 not n1308 ; n1308_not
g28757 not n4170 ; n4170_not
g28758 not n1281 ; n1281_not
g28759 not n1317 ; n1317_not
g28760 not n1065 ; n1065_not
g28761 not n1326 ; n1326_not
g28762 not n4161 ; n4161_not
g28763 not n1335 ; n1335_not
g28764 not n4152 ; n4152_not
g28765 not n4143 ; n4143_not
g28766 not n1353 ; n1353_not
g28767 not n3324 ; n3324_not
g28768 not n1029 ; n1029_not
g28769 not n3405 ; n3405_not
g28770 not n1803 ; n1803_not
g28771 not n1920 ; n1920_not
g28772 not n6114 ; n6114_not
g28773 not n3144 ; n3144_not
g28774 not n5421 ; n5421_not
g28775 not n3135 ; n3135_not
g28776 not n5412 ; n5412_not
g28777 not n5520 ; n5520_not
g28778 not n6321 ; n6321_not
g28779 not n3315 ; n3315_not
g28780 not n3423 ; n3423_not
g28781 not n1911 ; n1911_not
g28782 not n3126 ; n3126_not
g28783 not n9300 ; n9300_not
g28784 not n9111 ; n9111_not
g28785 not n7104 ; n7104_not
g28786 not n2028 ; n2028_not
g28787 not n6105 ; n6105_not
g28788 not n6411 ; n6411_not
g28789 not n6312 ; n6312_not
g28790 not n3351 ; n3351_not
g28791 not n3180 ; n3180_not
g28792 not n5430 ; n5430_not
g28793 not n1830 ; n1830_not
g28794 not n3360 ; n3360_not
g28795 not n3171 ; n3171_not
g28796 not n6303 ; n6303_not
g28797 not n8103 ; n8103_not
g28798 not n1821 ; n1821_not
g28799 not n5502 ; n5502_not
g28800 not n3162 ; n3162_not
g28801 not n5223 ; n5223_not
g28802 not n3333 ; n3333_not
g28803 not n6402 ; n6402_not
g28804 not n1812 ; n1812_not
g28805 not n9021 ; n9021_not
g28806 not n3216 ; n3216_not
g28807 not n3153 ; n3153_not
g28808 not n3234 ; n3234_not
g28809 not n3450 ; n3450_not
g28810 not n3108 ; n3108_not
g28811 not n8013 ; n8013_not
g28812 not n2073 ; n2073_not
g28813 not n6330 ; n6330_not
g28814 not n2082 ; n2082_not
g28815 not n9210 ; n9210_not
g28816 not n6420 ; n6420_not
g28817 not n8121 ; n8121_not
g28818 not n5007 ; n5007_not
g28819 not n8040 ; n8040_not
g28820 not n3252 ; n3252_not
g28821 not n2037 ; n2037_not
g28822 not n3432 ; n3432_not
g28823 not n5403 ; n5403_not
g28824 not n3225 ; n3225_not
g28825 not n9201 ; n9201_not
g28826 not n2046 ; n2046_not
g28827 not n1902 ; n1902_not
g28828 not n2055 ; n2055_not
g28829 not n3441 ; n3441_not
g28830 not n6313 ; n6313_not
g28831 not n5017 ; n5017_not
g28832 not n3190 ; n3190_not
g28833 not n2731 ; n2731_not
g28834 not n8212 ; n8212_not
g28835 not n4162 ; n4162_not
g28836 not n3055 ; n3055_not
g28837 not n4153 ; n4153_not
g28838 not n6205 ; n6205_not
g28839 not n3064 ; n3064_not
g28840 not n4063 ; n4063_not
g28841 not n5170 ; n5170_not
g28842 not n4108 ; n4108_not
g28843 not n2704 ; n2704_not
g28844 not n4117 ; n4117_not
g28845 not n4090 ; n4090_not
g28846 not n3235 ; n3235_not
g28847 not n2713 ; n2713_not
g28848 not n6322 ; n6322_not
g28849 not n3217 ; n3217_not
g28850 not n4135 ; n4135_not
g28851 not n4081 ; n4081_not
g28852 not n3244 ; n3244_not
g28853 not n8221 ; n8221_not
g28854 not n4540 ; n4540_not
g28855 not n6223 ; n6223_not
g28856 not n3208 ; n3208_not
g28857 not n6214 ; n6214_not
g28858 not n4144 ; n4144_not
g28859 not n4072 ; n4072_not
g28860 not n7024 ; n7024_not
g28861 not n7132 ; n7132_not
g28862 not n7060 ; n7060_not
g28863 not n7141 ; n7141_not
g28864 not n4261 ; n4261_not
g28865 not n4441 ; n4441_not
g28866 not n5242 ; n5242_not
g28867 not n8302 ; n8302_not
g28868 not n3109 ; n3109_not
g28869 not n4252 ; n4252_not
g28870 not n7042 ; n7042_not
g28871 not n5233 ; n5233_not
g28872 not n4243 ; n4243_not
g28873 not n3091 ; n3091_not
g28874 not n4315 ; n4315_not
g28875 not n5008 ; n5008_not
g28876 not n7033 ; n7033_not
g28877 not n4423 ; n4423_not
g28878 not n3082 ; n3082_not
g28879 not n2551 ; n2551_not
g28880 not n4306 ; n4306_not
g28881 not n8140 ; n8140_not
g28882 not n2560 ; n2560_not
g28883 not n5251 ; n5251_not
g28884 not n3073 ; n3073_not
g28885 not n7051 ; n7051_not
g28886 not n4207 ; n4207_not
g28887 not n3163 ; n3163_not
g28888 not n2641 ; n2641_not
g28889 not n4180 ; n4180_not
g28890 not n6304 ; n6304_not
g28891 not n4513 ; n4513_not
g28892 not n8005 ; n8005_not
g28893 not n2650 ; n2650_not
g28894 not n5215 ; n5215_not
g28895 not n3172 ; n3172_not
g28896 not n4351 ; n4351_not
g28897 not n4171 ; n4171_not
g28898 not n8131 ; n8131_not
g28899 not n5206 ; n5206_not
g28900 not n4522 ; n4522_not
g28901 not n4432 ; n4432_not
g28902 not n3127 ; n3127_not
g28903 not n2605 ; n2605_not
g28904 not n7114 ; n7114_not
g28905 not n4234 ; n4234_not
g28906 not n2614 ; n2614_not
g28907 not n4027 ; n4027_not
g28908 not n3145 ; n3145_not
g28909 not n4405 ; n4405_not
g28910 not n4225 ; n4225_not
g28911 not n3154 ; n3154_not
g28912 not n7150 ; n7150_not
g28913 not n4009 ; n4009_not
g28914 not n2434 ; n2434_not
g28915 not n2623 ; n2623_not
g28916 not n6403 ; n6403_not
g28917 not n2902 ; n2902_not
g28918 not n3523 ; n3523_not
g28919 not n3424 ; n3424_not
g28920 not n4603 ; n4603_not
g28921 not n3721 ; n3721_not
g28922 not n2911 ; n2911_not
g28923 not n2920 ; n2920_not
g28924 not n7600 ; n7600_not
g28925 not n5062 ; n5062_not
g28926 not n3703 ; n3703_not
g28927 not n6610 ; n6610_not
g28928 not n6601 ; n6601_not
g28929 not n6412 ; n6412_not
g28930 not n5053 ; n5053_not
g28931 not n8230 ; n8230_not
g28932 not n3820 ; n3820_not
g28933 not n4414 ; n4414_not
g28934 not n3361 ; n3361_not
g28935 not n3802 ; n3802_not
g28936 not n8122 ; n8122_not
g28937 not n3406 ; n3406_not
g28938 not n7501 ; n7501_not
g28939 not n7411 ; n7411_not
g28940 not n7510 ; n7510_not
g28941 not n4702 ; n4702_not
g28942 not n3541 ; n3541_not
g28943 not n8311 ; n8311_not
g28944 not n4711 ; n4711_not
g28945 not n6700 ; n6700_not
g28946 not n3433 ; n3433_not
g28947 not n4720 ; n4720_not
g28948 not n4900 ; n4900_not
g28949 not n6232 ; n6232_not
g28950 not n3460 ; n3460_not
g28951 not n8041 ; n8041_not
g28952 not n8203 ; n8203_not
g28953 not n3532 ; n3532_not
g28954 not n8032 ; n8032_not
g28955 not n8014 ; n8014_not
g28956 not n3505 ; n3505_not
g28957 not n3514 ; n3514_not
g28958 not n6430 ; n6430_not
g28959 not n3604 ; n3604_not
g28960 not n3442 ; n3442_not
g28961 not n4801 ; n4801_not
g28962 not n4810 ; n4810_not
g28963 not n3631 ; n3631_not
g28964 not n5026 ; n5026_not
g28965 not n5044 ; n5044_not
g28966 not n3613 ; n3613_not
g28967 not n8050 ; n8050_not
g28968 not n3451 ; n3451_not
g28969 not n6520 ; n6520_not
g28970 not n6511 ; n6511_not
g28971 not n6502 ; n6502_not
g28972 not n3226 ; n3226_not
g28973 not n8113 ; n8113_not
g28974 not n7213 ; n7213_not
g28975 not n5134 ; n5134_not
g28976 not n4450 ; n4450_not
g28977 not n6241 ; n6241_not
g28978 not n3037 ; n3037_not
g28979 not n7222 ; n7222_not
g28980 not n3307 ; n3307_not
g28981 not n2803 ; n2803_not
g28982 not n7231 ; n7231_not
g28983 not n8410 ; n8410_not
g28984 not n5125 ; n5125_not
g28985 not n3316 ; n3316_not
g28986 not n7123 ; n7123_not
g28987 not n2812 ; n2812_not
g28988 not n4054 ; n4054_not
g28989 not n7204 ; n7204_not
g28990 not n3253 ; n3253_not
g28991 not n3262 ; n3262_not
g28992 not n4036 ; n4036_not
g28993 not n8500 ; n8500_not
g28994 not n3046 ; n3046_not
g28995 not n5152 ; n5152_not
g28996 not n3271 ; n3271_not
g28997 not n3811 ; n3811_not
g28998 not n4018 ; n4018_not
g28999 not n4360 ; n4360_not
g29000 not n6331 ; n6331_not
g29001 not n3901 ; n3901_not
g29002 not n3352 ; n3352_not
g29003 not n3019 ; n3019_not
g29004 not n4612 ; n4612_not
g29005 not n5107 ; n5107_not
g29006 not n4621 ; n4621_not
g29007 not n4504 ; n4504_not
g29008 not n8104 ; n8104_not
g29009 not n4630 ; n4630_not
g29010 not n7402 ; n7402_not
g29011 not n3370 ; n3370_not
g29012 not n7420 ; n7420_not
g29013 not n7240 ; n7240_not
g29014 not n7015 ; n7015_not
g29015 not n3334 ; n3334_not
g29016 not n7006 ; n7006_not
g29017 not n8401 ; n8401_not
g29018 not n3028 ; n3028_not
g29019 not n2821 ; n2821_not
g29020 not n3325 ; n3325_not
g29021 not n5116 ; n5116_not
g29022 not n3343 ; n3343_not
g29023 not n7303 ; n7303_not
g29024 not n3910 ; n3910_not
g29025 not n7312 ; n7312_not
g29026 not n7321 ; n7321_not
g29027 not n1453 ; n1453_not
g29028 not n2281 ; n2281_not
g29029 not n1471 ; n1471_not
g29030 not n2326 ; n2326_not
g29031 not n1444 ; n1444_not
g29032 not n9202 ; n9202_not
g29033 not n1480 ; n1480_not
g29034 not n9211 ; n9211_not
g29035 not n5620 ; n5620_not
g29036 not n1507 ; n1507_not
g29037 not n1516 ; n1516_not
g29038 not n1534 ; n1534_not
g29039 not n1525 ; n1525_not
g29040 not n6106 ; n6106_not
g29041 not n9220 ; n9220_not
g29042 not n5611 ; n5611_not
g29043 not n1543 ; n1543_not
g29044 not n2254 ; n2254_not
g29045 not n2416 ; n2416_not
g29046 not n1462 ; n1462_not
g29047 not n1552 ; n1552_not
g29048 not n1354 ; n1354_not
g29049 not n1561 ; n1561_not
g29050 not n9031 ; n9031_not
g29051 not n1570 ; n1570_not
g29052 not n1840 ; n1840_not
g29053 not n1831 ; n1831_not
g29054 not n1255 ; n1255_not
g29055 not n1336 ; n1336_not
g29056 not n2461 ; n2461_not
g29057 not n1345 ; n1345_not
g29058 not n2272 ; n2272_not
g29059 not n2452 ; n2452_not
g29060 not n1372 ; n1372_not
g29061 not n1930 ; n1930_not
g29062 not n1381 ; n1381_not
g29063 not n5440 ; n5440_not
g29064 not n9040 ; n9040_not
g29065 not n1318 ; n1318_not
g29066 not n1417 ; n1417_not
g29067 not n1921 ; n1921_not
g29068 not n6043 ; n6043_not
g29069 not n6115 ; n6115_not
g29070 not n1903 ; n1903_not
g29071 not n1426 ; n1426_not
g29072 not n1435 ; n1435_not
g29073 not n1912 ; n1912_not
g29074 not n5323 ; n5323_not
g29075 not n1363 ; n1363_not
g29076 not n2443 ; n2443_not
g29077 not n9301 ; n9301_not
g29078 not n2380 ; n2380_not
g29079 not n9112 ; n9112_not
g29080 not n5521 ; n5521_not
g29081 not n2155 ; n2155_not
g29082 not n9400 ; n9400_not
g29083 not n6160 ; n6160_not
g29084 not n2317 ; n2317_not
g29085 not n2371 ; n2371_not
g29086 not n6052 ; n6052_not
g29087 not n5341 ; n5341_not
g29088 not n6070 ; n6070_not
g29089 not n2335 ; n2335_not
g29090 not n1705 ; n1705_not
g29091 not n1714 ; n1714_not
g29092 not n5530 ; n5530_not
g29093 not n6061 ; n6061_not
g29094 not n1732 ; n1732_not
g29095 not n1741 ; n1741_not
g29096 not n5305 ; n5305_not
g29097 not n2353 ; n2353_not
g29098 not n2245 ; n2245_not
g29099 not n5260 ; n5260_not
g29100 not n2290 ; n2290_not
g29101 not n6016 ; n6016_not
g29102 not n1723 ; n1723_not
g29103 not n2407 ; n2407_not
g29104 not n1615 ; n1615_not
g29105 not n1624 ; n1624_not
g29106 not n1822 ; n1822_not
g29107 not n1633 ; n1633_not
g29108 not n6151 ; n6151_not
g29109 not n5503 ; n5503_not
g29110 not n1606 ; n1606_not
g29111 not n9022 ; n9022_not
g29112 not n9004 ; n9004_not
g29113 not n1642 ; n1642_not
g29114 not n1813 ; n1813_not
g29115 not n1804 ; n1804_not
g29116 not n5512 ; n5512_not
g29117 not n6034 ; n6034_not
g29118 not n1660 ; n1660_not
g29119 not n5332 ; n5332_not
g29120 not n2362 ; n2362_not
g29121 not n2308 ; n2308_not
g29122 not n2056 ; n2056_not
g29123 not n2047 ; n2047_not
g29124 not n5404 ; n5404_not
g29125 not n1192 ; n1192_not
g29126 not n2029 ; n2029_not
g29127 not n5701 ; n5701_not
g29128 not n5800 ; n5800_not
g29129 not n1048 ; n1048_not
g29130 not n6007 ; n6007_not
g29131 not n1138 ; n1138_not
g29132 not n1039 ; n1039_not
g29133 not n6142 ; n6142_not
g29134 not n1219 ; n1219_not
g29135 not n1228 ; n1228_not
g29136 not n2182 ; n2182_not
g29137 not n2092 ; n2092_not
g29138 not n1129 ; n1129_not
g29139 not n2128 ; n2128_not
g29140 not n1246 ; n1246_not
g29141 not n9103 ; n9103_not
g29142 not n1084 ; n1084_not
g29143 not n2209 ; n2209_not
g29144 not n2515 ; n2515_not
g29145 not n2083 ; n2083_not
g29146 not n2218 ; n2218_not
g29147 not n2506 ; n2506_not
g29148 not n6124 ; n6124_not
g29149 not n1147 ; n1147_not
g29150 not n2074 ; n2074_not
g29151 not n1156 ; n1156_not
g29152 not n2227 ; n2227_not
g29153 not n1075 ; n1075_not
g29154 not n2038 ; n2038_not
g29155 not n1066 ; n1066_not
g29156 not n2236 ; n2236_not
g29157 not n2191 ; n2191_not
g29158 not n2065 ; n2065_not
g29159 not n1174 ; n1174_not
g29160 not n2524 ; n2524_not
g29161 not n1057 ; n1057_not
g29162 not n2470 ; n2470_not
g29163 not n2542 ; n2542_not
g29164 not n1282 ; n1282_not
g29165 not n5314 ; n5314_not
g29166 not n9121 ; n9121_not
g29167 not n1291 ; n1291_not
g29168 not n5224 ; n5224_not
g29169 not n5422 ; n5422_not
g29170 not n1309 ; n1309_not
g29171 not n2263 ; n2263_not
g29172 not n9130 ; n9130_not
g29173 not n2164 ; n2164_not
g29174 not n1327 ; n1327_not
g29175 not n2533 ; n2533_not
g29176 not n1264 ; n1264_not
g29177 not n6133 ; n6133_not
g29178 not n5413 ; n5413_not
g29179 not n2146 ; n2146_not
g29180 not n6413 ; n6413_not
g29181 not n2129 ; n2129_not
g29182 not n5531 ; n5531_not
g29183 not n8051 ; n8051_not
g29184 not n6134 ; n6134_not
g29185 not n4901 ; n4901_not
g29186 not n4721 ; n4721_not
g29187 not n3056 ; n3056_not
g29188 not n1814 ; n1814_not
g29189 not n1643 ; n1643_not
g29190 not n6071 ; n6071_not
g29191 not n1805 ; n1805_not
g29192 not n8024 ; n8024_not
g29193 not n5009 ; n5009_not
g29194 not n8141 ; n8141_not
g29195 not n2156 ; n2156_not
g29196 not n5522 ; n5522_not
g29197 not n3371 ; n3371_not
g29198 not n3092 ; n3092_not
g29199 not n2084 ; n2084_not
g29200 not n2165 ; n2165_not
g29201 not n3380 ; n3380_not
g29202 not n5504 ; n5504_not
g29203 not n3443 ; n3443_not
g29204 not n5540 ; n5540_not
g29205 not n3506 ; n3506_not
g29206 not n3434 ; n3434_not
g29207 not n9302 ; n9302_not
g29208 not n3470 ; n3470_not
g29209 not n6125 ; n6125_not
g29210 not n2093 ; n2093_not
g29211 not n9311 ; n9311_not
g29212 not n3461 ; n3461_not
g29213 not n6404 ; n6404_not
g29214 not n2147 ; n2147_not
g29215 not n1760 ; n1760_not
g29216 not n3083 ; n3083_not
g29217 not n3029 ; n3029_not
g29218 not n6152 ; n6152_not
g29219 not n9320 ; n9320_not
g29220 not n3425 ; n3425_not
g29221 not n2912 ; n2912_not
g29222 not n8033 ; n8033_not
g29223 not n3290 ; n3290_not
g29224 not n3416 ; n3416_not
g29225 not n6422 ; n6422_not
g29226 not n5513 ; n5513_not
g29227 not n3065 ; n3065_not
g29228 not n3452 ; n3452_not
g29229 not n3407 ; n3407_not
g29230 not n9122 ; n9122_not
g29231 not n1922 ; n1922_not
g29232 not n5414 ; n5414_not
g29233 not n1913 ; n1913_not
g29234 not n3128 ; n3128_not
g29235 not n3227 ; n3227_not
g29236 not n9113 ; n9113_not
g29237 not n1904 ; n1904_not
g29238 not n5450 ; n5450_not
g29239 not n9104 ; n9104_not
g29240 not n3236 ; n3236_not
g29241 not n6323 ; n6323_not
g29242 not n3119 ; n3119_not
g29243 not n3245 ; n3245_not
g29244 not n9203 ; n9203_not
g29245 not n5405 ; n5405_not
g29246 not n6314 ; n6314_not
g29247 not n9212 ; n9212_not
g29248 not n3254 ; n3254_not
g29249 not n8123 ; n8123_not
g29250 not n9140 ; n9140_not
g29251 not n6305 ; n6305_not
g29252 not n3173 ; n3173_not
g29253 not n3164 ; n3164_not
g29254 not n5432 ; n5432_not
g29255 not n8132 ; n8132_not
g29256 not n9131 ; n9131_not
g29257 not n4802 ; n4802_not
g29258 not n3191 ; n3191_not
g29259 not n1940 ; n1940_not
g29260 not n6116 ; n6116_not
g29261 not n3209 ; n3209_not
g29262 not n9032 ; n9032_not
g29263 not n5423 ; n5423_not
g29264 not n1931 ; n1931_not
g29265 not n3146 ; n3146_not
g29266 not n5441 ; n5441_not
g29267 not n3317 ; n3317_not
g29268 not n6044 ; n6044_not
g29269 not n5351 ; n5351_not
g29270 not n3326 ; n3326_not
g29271 not n2066 ; n2066_not
g29272 not n1841 ; n1841_not
g29273 not n1706 ; n1706_not
g29274 not n3335 ; n3335_not
g29275 not n1832 ; n1832_not
g29276 not n6350 ; n6350_not
g29277 not n2075 ; n2075_not
g29278 not n3353 ; n3353_not
g29279 not n3344 ; n3344_not
g29280 not n3362 ; n3362_not
g29281 not n1823 ; n1823_not
g29282 not n8105 ; n8105_not
g29283 not n6080 ; n6080_not
g29284 not n3263 ; n3263_not
g29285 not n6107 ; n6107_not
g29286 not n3272 ; n3272_not
g29287 not n6332 ; n6332_not
g29288 not n3281 ; n3281_not
g29289 not n8114 ; n8114_not
g29290 not n9221 ; n9221_not
g29291 not n2057 ; n2057_not
g29292 not n2921 ; n2921_not
g29293 not n9230 ; n9230_not
g29294 not n2039 ; n2039_not
g29295 not n1715 ; n1715_not
g29296 not n3308 ; n3308_not
g29297 not n1850 ; n1850_not
g29298 not n1346 ; n1346_not
g29299 not n4145 ; n4145_not
g29300 not n1337 ; n1337_not
g29301 not n4307 ; n4307_not
g29302 not n4523 ; n4523_not
g29303 not n1256 ; n1256_not
g29304 not n1328 ; n1328_not
g29305 not n4163 ; n4163_not
g29306 not n1319 ; n1319_not
g29307 not n1292 ; n1292_not
g29308 not n4514 ; n4514_not
g29309 not n1175 ; n1175_not
g29310 not n4181 ; n4181_not
g29311 not n4505 ; n4505_not
g29312 not n4370 ; n4370_not
g29313 not n4190 ; n4190_not
g29314 not n1283 ; n1283_not
g29315 not n7151 ; n7151_not
g29316 not n4208 ; n4208_not
g29317 not n5810 ; n5810_not
g29318 not n1274 ; n1274_not
g29319 not n4217 ; n4217_not
g29320 not n1265 ; n1265_not
g29321 not n4226 ; n4226_not
g29322 not n1463 ; n1463_not
g29323 not n4037 ; n4037_not
g29324 not n1454 ; n1454_not
g29325 not n4055 ; n4055_not
g29326 not n1445 ; n1445_not
g29327 not n7205 ; n7205_not
g29328 not n4073 ; n4073_not
g29329 not n1436 ; n1436_not
g29330 not n4541 ; n4541_not
g29331 not n4082 ; n4082_not
g29332 not n4064 ; n4064_not
g29333 not n7025 ; n7025_not
g29334 not n4091 ; n4091_not
g29335 not n9500 ; n9500_not
g29336 not n1382 ; n1382_not
g29337 not n4118 ; n4118_not
g29338 not n4109 ; n4109_not
g29339 not n1373 ; n1373_not
g29340 not n3911 ; n3911_not
g29341 not n1364 ; n1364_not
g29342 not n4127 ; n4127_not
g29343 not n4136 ; n4136_not
g29344 not n1355 ; n1355_not
g29345 not n5630 ; n5630_not
g29346 not n5900 ; n5900_not
g29347 not n1067 ; n1067_not
g29348 not n4352 ; n4352_not
g29349 not n1058 ; n1058_not
g29350 not n7061 ; n7061_not
g29351 not n1049 ; n1049_not
g29352 not n4361 ; n4361_not
g29353 not n5720 ; n5720_not
g29354 not n7016 ; n7016_not
g29355 not n4442 ; n4442_not
g29356 not n3641 ; n3641_not
g29357 not n7070 ; n7070_not
g29358 not n4433 ; n4433_not
g29359 not n2813 ; n2813_not
g29360 not n4406 ; n4406_not
g29361 not n4415 ; n4415_not
g29362 not n4424 ; n4424_not
g29363 not n1247 ; n1247_not
g29364 not n1238 ; n1238_not
g29365 not n5801 ; n5801_not
g29366 not n7043 ; n7043_not
g29367 not n5702 ; n5702_not
g29368 not n4262 ; n4262_not
g29369 not n7133 ; n7133_not
g29370 not n4280 ; n4280_not
g29371 not n5711 ; n5711_not
g29372 not n1157 ; n1157_not
g29373 not n4253 ; n4253_not
g29374 not n1148 ; n1148_not
g29375 not n1139 ; n1139_not
g29376 not n4316 ; n4316_not
g29377 not n4325 ; n4325_not
g29378 not n4460 ; n4460_not
g29379 not n1094 ; n1094_not
g29380 not n1085 ; n1085_not
g29381 not n4334 ; n4334_not
g29382 not n7115 ; n7115_not
g29383 not n1076 ; n1076_not
g29384 not n4451 ; n4451_not
g29385 not n3650 ; n3650_not
g29386 not n1670 ; n1670_not
g29387 not n7700 ; n7700_not
g29388 not n6602 ; n6602_not
g29389 not n6611 ; n6611_not
g29390 not n7610 ; n7610_not
g29391 not n6620 ; n6620_not
g29392 not n7601 ; n7601_not
g29393 not n3704 ; n3704_not
g29394 not n1661 ; n1661_not
g29395 not n3713 ; n3713_not
g29396 not n9410 ; n9410_not
g29397 not n6035 ; n6035_not
g29398 not n3722 ; n3722_not
g29399 not n1652 ; n1652_not
g29400 not n4730 ; n4730_not
g29401 not n3740 ; n3740_not
g29402 not n6701 ; n6701_not
g29403 not n7520 ; n7520_not
g29404 not n4703 ; n4703_not
g29405 not n6710 ; n6710_not
g29406 not n7511 ; n7511_not
g29407 not n7502 ; n7502_not
g29408 not n7412 ; n7412_not
g29409 not n6521 ; n6521_not
g29410 not n1634 ; n1634_not
g29411 not n1742 ; n1742_not
g29412 not n6431 ; n6431_not
g29413 not n1733 ; n1733_not
g29414 not n3524 ; n3524_not
g29415 not n6440 ; n6440_not
g29416 not n1724 ; n1724_not
g29417 not n6053 ; n6053_not
g29418 not n3542 ; n3542_not
g29419 not n8006 ; n8006_not
g29420 not n3560 ; n3560_not
g29421 not n6215 ; n6215_not
g29422 not n1562 ; n1562_not
g29423 not n6512 ; n6512_not
g29424 not n4820 ; n4820_not
g29425 not n6530 ; n6530_not
g29426 not n3605 ; n3605_not
g29427 not n3614 ; n3614_not
g29428 not n3623 ; n3623_not
g29429 not n4811 ; n4811_not
g29430 not n3632 ; n3632_not
g29431 not n1544 ; n1544_not
g29432 not n7304 ; n7304_not
g29433 not n1553 ; n1553_not
g29434 not n7007 ; n7007_not
g29435 not n5612 ; n5612_not
g29436 not n7241 ; n7241_not
g29437 not n1535 ; n1535_not
g29438 not n7124 ; n7124_not
g29439 not n7232 ; n7232_not
g29440 not n1526 ; n1526_not
g29441 not n7223 ; n7223_not
g29442 not n3812 ; n3812_not
g29443 not n7214 ; n7214_not
g29444 not n1517 ; n1517_not
g29445 not n4019 ; n4019_not
g29446 not n1481 ; n1481_not
g29447 not n1472 ; n1472_not
g29448 not n4028 ; n4028_not
g29449 not n3803 ; n3803_not
g29450 not n6800 ; n6800_not
g29451 not n6026 ; n6026_not
g29452 not n1625 ; n1625_not
g29453 not n3821 ; n3821_not
g29454 not n7421 ; n7421_not
g29455 not n1616 ; n1616_not
g29456 not n1607 ; n1607_not
g29457 not n4640 ; n4640_not
g29458 not n4631 ; n4631_not
g29459 not n6017 ; n6017_not
g29460 not n4622 ; n4622_not
g29461 not n4613 ; n4613_not
g29462 not n7340 ; n7340_not
g29463 not n7331 ; n7331_not
g29464 not n7322 ; n7322_not
g29465 not n3902 ; n3902_not
g29466 not n4604 ; n4604_not
g29467 not n1571 ; n1571_not
g29468 not n7313 ; n7313_not
g29469 not n3920 ; n3920_not
g29470 not n2624 ; n2624_not
g29471 not n5225 ; n5225_not
g29472 not n5144 ; n5144_not
g29473 not n5315 ; n5315_not
g29474 not n5045 ; n5045_not
g29475 not n2462 ; n2462_not
g29476 not n8312 ; n8312_not
g29477 not n2642 ; n2642_not
g29478 not n9023 ; n9023_not
g29479 not n8222 ; n8222_not
g29480 not n2453 ; n2453_not
g29481 not n5162 ; n5162_not
g29482 not n6008 ; n6008_not
g29483 not n8231 ; n8231_not
g29484 not n8150 ; n8150_not
g29485 not n5090 ; n5090_not
g29486 not n5360 ; n5360_not
g29487 not n5207 ; n5207_not
g29488 not n6161 ; n6161_not
g29489 not n5153 ; n5153_not
g29490 not n2228 ; n2228_not
g29491 not n2318 ; n2318_not
g29492 not n2255 ; n2255_not
g29493 not n6170 ; n6170_not
g29494 not n5234 ; n5234_not
g29495 not n8420 ; n8420_not
g29496 not n2606 ; n2606_not
g29497 not n2264 ; n2264_not
g29498 not n8213 ; n8213_not
g29499 not n8330 ; n8330_not
g29500 not n2309 ; n2309_not
g29501 not n2480 ; n2480_not
g29502 not n2381 ; n2381_not
g29503 not n2615 ; n2615_not
g29504 not n5306 ; n5306_not
g29505 not n2471 ; n2471_not
g29506 not n5135 ; n5135_not
g29507 not n9005 ; n9005_not
g29508 not n8321 ; n8321_not
g29509 not n5063 ; n5063_not
g29510 not n2390 ; n2390_not
g29511 not n2750 ; n2750_not
g29512 not n5180 ; n5180_not
g29513 not n2930 ; n2930_not
g29514 not n2291 ; n2291_not
g29515 not n2417 ; n2417_not
g29516 not n2714 ; n2714_not
g29517 not n2741 ; n2741_not
g29518 not n5171 ; n5171_not
g29519 not n2723 ; n2723_not
g29520 not n6224 ; n6224_not
g29521 not n5072 ; n5072_not
g29522 not n2408 ; n2408_not
g29523 not n8510 ; n8510_not
g29524 not n5261 ; n5261_not
g29525 not n2732 ; n2732_not
g29526 not n6260 ; n6260_not
g29527 not n5054 ; n5054_not
g29528 not n8303 ; n8303_not
g29529 not n6233 ; n6233_not
g29530 not n8015 ; n8015_not
g29531 not n8240 ; n8240_not
g29532 not n8600 ; n8600_not
g29533 not n5324 ; n5324_not
g29534 not n2903 ; n2903_not
g29535 not n2444 ; n2444_not
g29536 not n2561 ; n2561_not
g29537 not n6206 ; n6206_not
g29538 not n2282 ; n2282_not
g29539 not n2435 ; n2435_not
g29540 not n2327 ; n2327_not
g29541 not n2705 ; n2705_not
g29542 not n5081 ; n5081_not
g29543 not n2570 ; n2570_not
g29544 not n9041 ; n9041_not
g29545 not n5342 ; n5342_not
g29546 not n6143 ; n6143_not
g29547 not n2219 ; n2219_not
g29548 not n2336 ; n2336_not
g29549 not n2363 ; n2363_not
g29550 not n5108 ; n5108_not
g29551 not n2237 ; n2237_not
g29552 not n2507 ; n2507_not
g29553 not n5027 ; n5027_not
g29554 not n5243 ; n5243_not
g29555 not n5126 ; n5126_not
g29556 not n3047 ; n3047_not
g29557 not n2840 ; n2840_not
g29558 not n5117 ; n5117_not
g29559 not n6242 ; n6242_not
g29560 not n2543 ; n2543_not
g29561 not n2354 ; n2354_not
g29562 not n5270 ; n5270_not
g29563 not n3038 ; n3038_not
g29564 not n2345 ; n2345_not
g29565 not n2525 ; n2525_not
g29566 not n2552 ; n2552_not
g29567 not n2822 ; n2822_not
g29568 not n2183 ; n2183_not
g29569 not n2516 ; n2516_not
g29570 not n5333 ; n5333_not
g29571 not n2246 ; n2246_not
g29572 not n8042 ; n8042_not
g29573 not n5036 ; n5036_not
g29574 not n2372 ; n2372_not
g29575 not n2804 ; n2804_not
g29576 not n2192 ; n2192_not
g29577 not n9006 ; n9006_not
g29578 not n3651 ; n3651_not
g29579 not n6810 ; n6810_not
g29580 not n3831 ; n3831_not
g29581 not n7422 ; n7422_not
g29582 not n1716 ; n1716_not
g29583 not n3543 ; n3543_not
g29584 not n6162 ; n6162_not
g29585 not n3642 ; n3642_not
g29586 not n2823 ; n2823_not
g29587 not n6531 ; n6531_not
g29588 not n7413 ; n7413_not
g29589 not n4641 ; n4641_not
g29590 not n6054 ; n6054_not
g29591 not n3804 ; n3804_not
g29592 not n7701 ; n7701_not
g29593 not n7152 ; n7152_not
g29594 not n3624 ; n3624_not
g29595 not n6351 ; n6351_not
g29596 not n1626 ; n1626_not
g29597 not n3615 ; n3615_not
g29598 not n2652 ; n2652_not
g29599 not n6234 ; n6234_not
g29600 not n6540 ; n6540_not
g29601 not n7440 ; n7440_not
g29602 not n3552 ; n3552_not
g29603 not n3813 ; n3813_not
g29604 not n8304 ; n8304_not
g29605 not n4803 ; n4803_not
g29606 not n3822 ; n3822_not
g29607 not n4650 ; n4650_not
g29608 not n7431 ; n7431_not
g29609 not n8007 ; n8007_not
g29610 not n4614 ; n4614_not
g29611 not n5172 ; n5172_not
g29612 not n7053 ; n7053_not
g29613 not n2832 ; n2832_not
g29614 not n6009 ; n6009_not
g29615 not n5118 ; n5118_not
g29616 not n5802 ; n5802_not
g29617 not n7341 ; n7341_not
g29618 not n4812 ; n4812_not
g29619 not n8106 ; n8106_not
g29620 not n1743 ; n1743_not
g29621 not n1581 ; n1581_not
g29622 not n8511 ; n8511_not
g29623 not n7332 ; n7332_not
g29624 not n4515 ; n4515_not
g29625 not n3660 ; n3660_not
g29626 not n3507 ; n3507_not
g29627 not n7323 ; n7323_not
g29628 not n2409 ; n2409_not
g29629 not n3318 ; n3318_not
g29630 not n5163 ; n5163_not
g29631 not n6450 ; n6450_not
g29632 not n1608 ; n1608_not
g29633 not n6441 ; n6441_not
g29634 not n6018 ; n6018_not
g29635 not n2742 ; n2742_not
g29636 not n9303 ; n9303_not
g29637 not n3840 ; n3840_not
g29638 not n1725 ; n1725_not
g29639 not n4623 ; n4623_not
g29640 not n5127 ; n5127_not
g29641 not n8403 ; n8403_not
g29642 not n3525 ; n3525_not
g29643 not n1590 ; n1590_not
g29644 not n9015 ; n9015_not
g29645 not n5334 ; n5334_not
g29646 not n7350 ; n7350_not
g29647 not n9420 ; n9420_not
g29648 not n4830 ; n4830_not
g29649 not n2625 ; n2625_not
g29650 not n6513 ; n6513_not
g29651 not n6045 ; n6045_not
g29652 not n3390 ; n3390_not
g29653 not n3723 ; n3723_not
g29654 not n4605 ; n4605_not
g29655 not n3732 ; n3732_not
g29656 not n2364 ; n2364_not
g29657 not n5145 ; n5145_not
g29658 not n4731 ; n4731_not
g29659 not n4722 ; n4722_not
g29660 not n1653 ; n1653_not
g29661 not n6603 ; n6603_not
g29662 not n1671 ; n1671_not
g29663 not n5550 ; n5550_not
g29664 not n9123 ; n9123_not
g29665 not n3741 ; n3741_not
g29666 not n6504 ; n6504_not
g29667 not n7611 ; n7611_not
g29668 not n7620 ; n7620_not
g29669 not n2382 ; n2382_not
g29670 not n3480 ; n3480_not
g29671 not n6630 ; n6630_not
g29672 not n7602 ; n7602_not
g29673 not n9411 ; n9411_not
g29674 not n1662 ; n1662_not
g29675 not n3606 ; n3606_not
g29676 not n6612 ; n6612_not
g29677 not n8133 ; n8133_not
g29678 not n3705 ; n3705_not
g29679 not n8430 ; n8430_not
g29680 not n6621 ; n6621_not
g29681 not n3273 ; n3273_not
g29682 not n3714 ; n3714_not
g29683 not n2814 ; n2814_not
g29684 not n6243 ; n6243_not
g29685 not n2481 ; n2481_not
g29686 not n4632 ; n4632_not
g29687 not n4452 ; n4452_not
g29688 not n9402 ; n9402_not
g29689 not n8421 ; n8421_not
g29690 not n6522 ; n6522_not
g29691 not n5154 ; n5154_not
g29692 not n4434 ; n4434_not
g29693 not n3561 ; n3561_not
g29694 not n1635 ; n1635_not
g29695 not n1680 ; n1680_not
g29696 not n5343 ; n5343_not
g29697 not n7710 ; n7710_not
g29698 not n2760 ; n2760_not
g29699 not n7233 ; n7233_not
g29700 not n7530 ; n7530_not
g29701 not n6702 ; n6702_not
g29702 not n6027 ; n6027_not
g29703 not n4704 ; n4704_not
g29704 not n1644 ; n1644_not
g29705 not n7512 ; n7512_not
g29706 not n9330 ; n9330_not
g29707 not n7215 ; n7215_not
g29708 not n6711 ; n6711_not
g29709 not n7125 ; n7125_not
g29710 not n2391 ; n2391_not
g29711 not n1617 ; n1617_not
g29712 not n7503 ; n7503_not
g29713 not n1707 ; n1707_not
g29714 not n3381 ; n3381_not
g29715 not n6720 ; n6720_not
g29716 not n2490 ; n2490_not
g29717 not n8700 ; n8700_not
g29718 not n1149 ; n1149_not
g29719 not n7035 ; n7035_not
g29720 not n1086 ; n1086_not
g29721 not n1194 ; n1194_not
g29722 not n7044 ; n7044_not
g29723 not n4254 ; n4254_not
g29724 not n6171 ; n6171_not
g29725 not n4263 ; n4263_not
g29726 not n4083 ; n4083_not
g29727 not n1185 ; n1185_not
g29728 not n4272 ; n4272_not
g29729 not n7134 ; n7134_not
g29730 not n4281 ; n4281_not
g29731 not n1176 ; n1176_not
g29732 not n1068 ; n1068_not
g29733 not n4236 ; n4236_not
g29734 not n4470 ; n4470_not
g29735 not n5244 ; n5244_not
g29736 not n4038 ; n4038_not
g29737 not n4506 ; n4506_not
g29738 not n5316 ; n5316_not
g29739 not n4191 ; n4191_not
g29740 not n2436 ; n2436_not
g29741 not n5811 ; n5811_not
g29742 not n1284 ; n1284_not
g29743 not n5307 ; n5307_not
g29744 not n4209 ; n4209_not
g29745 not n1275 ; n1275_not
g29746 not n2616 ; n2616_not
g29747 not n4218 ; n4218_not
g29748 not n1266 ; n1266_not
g29749 not n2454 ; n2454_not
g29750 not n2607 ; n2607_not
g29751 not n4227 ; n4227_not
g29752 not n1257 ; n1257_not
g29753 not n1239 ; n1239_not
g29754 not n2526 ; n2526_not
g29755 not n7107 ; n7107_not
g29756 not n2553 ; n2553_not
g29757 not n4371 ; n4371_not
g29758 not n4290 ; n4290_not
g29759 not n5451 ; n5451_not
g29760 not n4380 ; n4380_not
g29761 not n4443 ; n4443_not
g29762 not n5262 ; n5262_not
g29763 not n5181 ; n5181_not
g29764 not n5271 ; n5271_not
g29765 not n7080 ; n7080_not
g29766 not n2544 ; n2544_not
g29767 not n5055 ; n5055_not
g29768 not n4407 ; n4407_not
g29769 not n7071 ; n7071_not
g29770 not n2535 ; n2535_not
g29771 not n4416 ; n4416_not
g29772 not n1356 ; n1356_not
g29773 not n6180 ; n6180_not
g29774 not n4425 ; n4425_not
g29775 not n5712 ; n5712_not
g29776 not n1167 ; n1167_not
g29777 not n1158 ; n1158_not
g29778 not n4308 ; n4308_not
g29779 not n2580 ; n2580_not
g29780 not n4317 ; n4317_not
g29781 not n1095 ; n1095_not
g29782 not n4326 ; n4326_not
g29783 not n2508 ; n2508_not
g29784 not n4461 ; n4461_not
g29785 not n5721 ; n5721_not
g29786 not n2517 ; n2517_not
g29787 not n4335 ; n4335_not
g29788 not n1077 ; n1077_not
g29789 not n2571 ; n2571_not
g29790 not n4344 ; n4344_not
g29791 not n7062 ; n7062_not
g29792 not n2562 ; n2562_not
g29793 not n4353 ; n4353_not
g29794 not n2418 ; n2418_not
g29795 not n7017 ; n7017_not
g29796 not n7242 ; n7242_not
g29797 not n1536 ; n1536_not
g29798 not n2427 ; n2427_not
g29799 not n1527 ; n1527_not
g29800 not n7224 ; n7224_not
g29801 not n5613 ; n5613_not
g29802 not n4551 ; n4551_not
g29803 not n2706 ; n2706_not
g29804 not n9213 ; n9213_not
g29805 not n9600 ; n9600_not
g29806 not n5703 ; n5703_not
g29807 not n1482 ; n1482_not
g29808 not n6216 ; n6216_not
g29809 not n5631 ; n5631_not
g29810 not n5190 ; n5190_not
g29811 not n4029 ; n4029_not
g29812 not n1464 ; n1464_not
g29813 not n9510 ; n9510_not
g29814 not n4920 ; n4920_not
g29815 not n3903 ; n3903_not
g29816 not n2733 ; n2733_not
g29817 not n1572 ; n1572_not
g29818 not n7314 ; n7314_not
g29819 not n3912 ; n3912_not
g29820 not n5604 ; n5604_not
g29821 not n3921 ; n3921_not
g29822 not n6225 ; n6225_not
g29823 not n6900 ; n6900_not
g29824 not n7305 ; n7305_not
g29825 not n6207 ; n6207_not
g29826 not n1563 ; n1563_not
g29827 not n2724 ; n2724_not
g29828 not n5910 ; n5910_not
g29829 not n1473 ; n1473_not
g29830 not n7008 ; n7008_not
g29831 not n1545 ; n1545_not
g29832 not n7260 ; n7260_not
g29833 not n4560 ; n4560_not
g29834 not n5370 ; n5370_not
g29835 not n1383 ; n1383_not
g29836 not n4119 ; n4119_not
g29837 not n2643 ; n2643_not
g29838 not n8610 ; n8610_not
g29839 not n1365 ; n1365_not
g29840 not n4128 ; n4128_not
g29841 not n5901 ; n5901_not
g29842 not n1347 ; n1347_not
g29843 not n1338 ; n1338_not
g29844 not n4146 ; n4146_not
g29845 not n2463 ; n2463_not
g29846 not n1329 ; n1329_not
g29847 not n4524 ; n4524_not
g29848 not n5226 ; n5226_not
g29849 not n2634 ; n2634_not
g29850 not n4164 ; n4164_not
g29851 not n1293 ; n1293_not
g29852 not n4182 ; n4182_not
g29853 not n5640 ; n5640_not
g29854 not n1455 ; n1455_not
g29855 not n4047 ; n4047_not
g29856 not n7206 ; n7206_not
g29857 not n4056 ; n4056_not
g29858 not n1374 ; n1374_not
g29859 not n1446 ; n1446_not
g29860 not n2445 ; n2445_not
g29861 not n4065 ; n4065_not
g29862 not n4542 ; n4542_not
g29863 not n1437 ; n1437_not
g29864 not n8601 ; n8601_not
g29865 not n4074 ; n4074_not
g29866 not n2670 ; n2670_not
g29867 not n1419 ; n1419_not
g29868 not n5208 ; n5208_not
g29869 not n4533 ; n4533_not
g29870 not n5730 ; n5730_not
g29871 not n4092 ; n4092_not
g29872 not n1392 ; n1392_not
g29873 not n8115 ; n8115_not
g29874 not n5064 ; n5064_not
g29875 not n3291 ; n3291_not
g29876 not n3237 ; n3237_not
g29877 not n5415 ; n5415_not
g29878 not n1824 ; n1824_not
g29879 not n9231 ; n9231_not
g29880 not n3309 ; n3309_not
g29881 not n5073 ; n5073_not
g29882 not n1851 ; n1851_not
g29883 not n2922 ; n2922_not
g29884 not n9240 ; n9240_not
g29885 not n3327 ; n3327_not
g29886 not n1842 ; n1842_not
g29887 not n6261 ; n6261_not
g29888 not n3336 ; n3336_not
g29889 not n1833 ; n1833_not
g29890 not n2913 ; n2913_not
g29891 not n5820 ; n5820_not
g29892 not n3066 ; n3066_not
g29893 not n6324 ; n6324_not
g29894 not n9204 ; n9204_not
g29895 not n6117 ; n6117_not
g29896 not n3255 ; n3255_not
g29897 not n2940 ; n2940_not
g29898 not n8250 ; n8250_not
g29899 not n3264 ; n3264_not
g29900 not n5460 ; n5460_not
g29901 not n6108 ; n6108_not
g29902 not n2283 ; n2283_not
g29903 not n6333 ; n6333_not
g29904 not n2931 ; n2931_not
g29905 not n3282 ; n3282_not
g29906 not n6342 ; n6342_not
g29907 not n5505 ; n5505_not
g29908 not n1806 ; n1806_not
g29909 not n8313 ; n8313_not
g29910 not n5091 ; n5091_not
g29911 not n3408 ; n3408_not
g29912 not n4911 ; n4911_not
g29913 not n8061 ; n8061_not
g29914 not n8322 ; n8322_not
g29915 not n3417 ; n3417_not
g29916 not n6405 ; n6405_not
g29917 not n9132 ; n9132_not
g29918 not n8052 ; n8052_not
g29919 not n8331 ; n8331_not
g29920 not n3435 ; n3435_not
g29921 not n6252 ; n6252_not
g29922 not n8340 ; n8340_not
g29923 not n3345 ; n3345_not
g29924 not n5082 ; n5082_not
g29925 not n3354 ; n3354_not
g29926 not n4902 ; n4902_not
g29927 not n6081 ; n6081_not
g29928 not n6360 ; n6360_not
g29929 not n1734 ; n1734_not
g29930 not n5352 ; n5352_not
g29931 not n8016 ; n8016_not
g29932 not n2715 ; n2715_not
g29933 not n3372 ; n3372_not
g29934 not n1815 ; n1815_not
g29935 not n9024 ; n9024_not
g29936 not n8070 ; n8070_not
g29937 not n2058 ; n2058_not
g29938 not n2067 ; n2067_not
g29939 not n2229 ; n2229_not
g29940 not n2238 ; n2238_not
g29941 not n8160 ; n8160_not
g29942 not n2049 ; n2049_not
g29943 not n5028 ; n5028_not
g29944 not n2193 ; n2193_not
g29945 not n5406 ; n5406_not
g29946 not n2247 ; n2247_not
g29947 not n9105 ; n9105_not
g29948 not n5136 ; n5136_not
g29949 not n3129 ; n3129_not
g29950 not n3138 ; n3138_not
g29951 not n2256 ; n2256_not
g29952 not n3048 ; n3048_not
g29953 not n2166 ; n2166_not
g29954 not n2175 ; n2175_not
g29955 not n9051 ; n9051_not
g29956 not n3057 ; n3057_not
g29957 not n2148 ; n2148_not
g29958 not n8151 ; n8151_not
g29959 not n2139 ; n2139_not
g29960 not n3039 ; n3039_not
g29961 not n9060 ; n9060_not
g29962 not n3075 ; n3075_not
g29963 not n2094 ; n2094_not
g29964 not n2184 ; n2184_not
g29965 not n3084 ; n3084_not
g29966 not n6126 ; n6126_not
g29967 not n9042 ; n9042_not
g29968 not n2085 ; n2085_not
g29969 not n5433 ; n5433_not
g29970 not n3183 ; n3183_not
g29971 not n9150 ; n9150_not
g29972 not n3192 ; n3192_not
g29973 not n5046 ; n5046_not
g29974 not n6315 ; n6315_not
g29975 not n1941 ; n1941_not
g29976 not n6135 ; n6135_not
g29977 not n1932 ; n1932_not
g29978 not n8223 ; n8223_not
g29979 not n5442 ; n5442_not
g29980 not n5361 ; n5361_not
g29981 not n1923 ; n1923_not
g29982 not n8232 ; n8232_not
g29983 not n1914 ; n1914_not
g29984 not n3228 ; n3228_not
g29985 not n1905 ; n1905_not
g29986 not n5235 ; n5235_not
g29987 not n9033 ; n9033_not
g29988 not n6144 ; n6144_not
g29989 not n3147 ; n3147_not
g29990 not n5424 ; n5424_not
g29991 not n8214 ; n8214_not
g29992 not n8043 ; n8043_not
g29993 not n3165 ; n3165_not
g29994 not n9141 ; n9141_not
g29995 not n1950 ; n1950_not
g29996 not n2265 ; n2265_not
g29997 not n3174 ; n3174_not
g29998 not n6306 ; n6306_not
g29999 not n6270 ; n6270_not
g30000 not n1752 ; n1752_not
g30001 not n3471 ; n3471_not
g30002 not n1770 ; n1770_not
g30003 not n9312 ; n9312_not
g30004 not n6153 ; n6153_not
g30005 not n8025 ; n8025_not
g30006 not n6423 ; n6423_not
g30007 not n2328 ; n2328_not
g30008 not n6414 ; n6414_not
g30009 not n5109 ; n5109_not
g30010 not n8034 ; n8034_not
g30011 not n2850 ; n2850_not
g30012 not n2346 ; n2346_not
g30013 not n3453 ; n3453_not
g30014 not n5523 ; n5523_not
g30015 not n2337 ; n2337_not
g30016 not n1761 ; n1761_not
g30017 not n5514 ; n5514_not
g30018 not n5532 ; n5532_not
g30019 not n9321 ; n9321_not
g30020 not n3462 ; n3462_not
g30021 not n1375 ; n1375_not
g30022 not n3049 ; n3049_not
g30023 not n9007 ; n9007_not
g30024 not n4066 ; n4066_not
g30025 not n5056 ; n5056_not
g30026 not n5911 ; n5911_not
g30027 not n2059 ; n2059_not
g30028 not n1096 ; n1096_not
g30029 not n3580 ; n3580_not
g30030 not n1438 ; n1438_not
g30031 not n1456 ; n1456_not
g30032 not n5920 ; n5920_not
g30033 not n2941 ; n2941_not
g30034 not n6109 ; n6109_not
g30035 not n6505 ; n6505_not
g30036 not n4048 ; n4048_not
g30037 not n5272 ; n5272_not
g30038 not n4327 ; n4327_not
g30039 not n5533 ; n5533_not
g30040 not n8242 ; n8242_not
g30041 not n6325 ; n6325_not
g30042 not n1564 ; n1564_not
g30043 not n8341 ; n8341_not
g30044 not n4543 ; n4543_not
g30045 not n1447 ; n1447_not
g30046 not n4318 ; n4318_not
g30047 not n4534 ; n4534_not
g30048 not n5650 ; n5650_not
g30049 not n6217 ; n6217_not
g30050 not n1915 ; n1915_not
g30051 not n2662 ; n2662_not
g30052 not n4093 ; n4093_not
g30053 not n8422 ; n8422_not
g30054 not n5641 ; n5641_not
g30055 not n9610 ; n9610_not
g30056 not n7180 ; n7180_not
g30057 not n5209 ; n5209_not
g30058 not n9016 ; n9016_not
g30059 not n9034 ; n9034_not
g30060 not n3571 ; n3571_not
g30061 not n9700 ; n9700_not
g30062 not n8404 ; n8404_not
g30063 not n1393 ; n1393_not
g30064 not n1384 ; n1384_not
g30065 not n5713 ; n5713_not
g30066 not n5452 ; n5452_not
g30067 not n8017 ; n8017_not
g30068 not n3472 ; n3472_not
g30069 not n2671 ; n2671_not
g30070 not n4840 ; n4840_not
g30071 not n2581 ; n2581_not
g30072 not n7126 ; n7126_not
g30073 not n1429 ; n1429_not
g30074 not n8602 ; n8602_not
g30075 not n1906 ; n1906_not
g30076 not n8224 ; n8224_not
g30077 not n2950 ; n2950_not
g30078 not n4084 ; n4084_not
g30079 not n3229 ; n3229_not
g30080 not n3526 ; n3526_not
g30081 not n8233 ; n8233_not
g30082 not n7027 ; n7027_not
g30083 not n7234 ; n7234_not
g30084 not n7801 ; n7801_not
g30085 not n4345 ; n4345_not
g30086 not n4219 ; n4219_not
g30087 not n1528 ; n1528_not
g30088 not n3283 ; n3283_not
g30089 not n4552 ; n4552_not
g30090 not n2194 ; n2194_not
g30091 not n1519 ; n1519_not
g30092 not n7810 ; n7810_not
g30093 not n5326 ; n5326_not
g30094 not n4822 ; n4822_not
g30095 not n2086 ; n2086_not
g30096 not n2707 ; n2707_not
g30097 not n8107 ; n8107_not
g30098 not n3274 ; n3274_not
g30099 not n7216 ; n7216_not
g30100 not n2284 ; n2284_not
g30101 not n6514 ; n6514_not
g30102 not n3292 ; n3292_not
g30103 not n4453 ; n4453_not
g30104 not n4561 ; n4561_not
g30105 not n2815 ; n2815_not
g30106 not n5065 ; n5065_not
g30107 not n9070 ; n9070_not
g30108 not n3238 ; n3238_not
g30109 not n7252 ; n7252_not
g30110 not n1537 ; n1537_not
g30111 not n8116 ; n8116_not
g30112 not n7243 ; n7243_not
g30113 not n5551 ; n5551_not
g30114 not n2419 ; n2419_not
g30115 not n3823 ; n3823_not
g30116 not n7063 ; n7063_not
g30117 not n6334 ; n6334_not
g30118 not n7018 ; n7018_not
g30119 not n2428 ; n2428_not
g30120 not n5182 ; n5182_not
g30121 not n3094 ; n3094_not
g30122 not n8251 ; n8251_not
g30123 not n8530 ; n8530_not
g30124 not n6415 ; n6415_not
g30125 not n2437 ; n2437_not
g30126 not n2833 ; n2833_not
g30127 not n5632 ; n5632_not
g30128 not n5191 ; n5191_not
g30129 not n6307 ; n6307_not
g30130 not n8710 ; n8710_not
g30131 not n6208 ; n6208_not
g30132 not n8701 ; n8701_not
g30133 not n1087 ; n1087_not
g30134 not n1465 ; n1465_not
g30135 not n5092 ; n5092_not
g30136 not n3931 ; n3931_not
g30137 not n4462 ; n4462_not
g30138 not n2068 ; n2068_not
g30139 not n1816 ; n1816_not
g30140 not n4831 ; n4831_not
g30141 not n9214 ; n9214_not
g30142 not n5614 ; n5614_not
g30143 not n6064 ; n6064_not
g30144 not n1078 ; n1078_not
g30145 not n5722 ; n5722_not
g30146 not n3256 ; n3256_not
g30147 not n9601 ; n9601_not
g30148 not n5623 ; n5623_not
g30149 not n1069 ; n1069_not
g30150 not n5461 ; n5461_not
g30151 not n1492 ; n1492_not
g30152 not n3265 ; n3265_not
g30153 not n2572 ; n2572_not
g30154 not n1483 ; n1483_not
g30155 not n1951 ; n1951_not
g30156 not n1960 ; n1960_not
g30157 not n2590 ; n2590_not
g30158 not n7054 ; n7054_not
g30159 not n5425 ; n5425_not
g30160 not n9133 ; n9133_not
g30161 not n3553 ; n3553_not
g30162 not n5407 ; n5407_not
g30163 not n4228 ; n4228_not
g30164 not n6091 ; n6091_not
g30165 not n3157 ; n3157_not
g30166 not n1258 ; n1258_not
g30167 not n3409 ; n3409_not
g30168 not n2482 ; n2482_not
g30169 not n6145 ; n6145_not
g30170 not n2824 ; n2824_not
g30171 not n3148 ; n3148_not
g30172 not n9520 ; n9520_not
g30173 not n8026 ; n8026_not
g30174 not n4471 ; n4471_not
g30175 not n8134 ; n8134_not
g30176 not n8215 ; n8215_not
g30177 not n5803 ; n5803_not
g30178 not n1168 ; n1168_not
g30179 not n5812 ; n5812_not
g30180 not n9142 ; n9142_not
g30181 not n1861 ; n1861_not
g30182 not n6118 ; n6118_not
g30183 not n2617 ; n2617_not
g30184 not n1276 ; n1276_not
g30185 not n3535 ; n3535_not
g30186 not n6460 ; n6460_not
g30187 not n3166 ; n3166_not
g30188 not n2158 ; n2158_not
g30189 not n3139 ; n3139_not
g30190 not n1573 ; n1573_not
g30191 not n1186 ; n1186_not
g30192 not n5704 ; n5704_not
g30193 not n5416 ; n5416_not
g30194 not n5236 ; n5236_not
g30195 not n7045 ; n7045_not
g30196 not n8206 ; n8206_not
g30197 not n4273 ; n4273_not
g30198 not n9106 ; n9106_not
g30199 not n7135 ; n7135_not
g30200 not n1177 ; n1177_not
g30201 not n5371 ; n5371_not
g30202 not n9340 ; n9340_not
g30203 not n2248 ; n2248_not
g30204 not n9115 ; n9115_not
g30205 not n6424 ; n6424_not
g30206 not n6163 ; n6163_not
g30207 not n4237 ; n4237_not
g30208 not n8800 ; n8800_not
g30209 not n4183 ; n4183_not
g30210 not n6154 ; n6154_not
g30211 not n4291 ; n4291_not
g30212 not n8008 ; n8008_not
g30213 not n6451 ; n6451_not
g30214 not n4246 ; n4246_not
g30215 not n3490 ; n3490_not
g30216 not n2257 ; n2257_not
g30217 not n3544 ; n3544_not
g30218 not n1195 ; n1195_not
g30219 not n9124 ; n9124_not
g30220 not n5344 ; n5344_not
g30221 not n1717 ; n1717_not
g30222 not n4255 ; n4255_not
g30223 not n6442 ; n6442_not
g30224 not n7144 ; n7144_not
g30225 not n2473 ; n2473_not
g30226 not n5317 ; n5317_not
g30227 not n4309 ; n4309_not
g30228 not n8125 ; n8125_not
g30229 not n2491 ; n2491_not
g30230 not n2644 ; n2644_not
g30231 not n1339 ; n1339_not
g30232 not n2347 ; n2347_not
g30233 not n4147 ; n4147_not
g30234 not n5245 ; n5245_not
g30235 not n6316 ; n6316_not
g30236 not n1726 ; n1726_not
g30237 not n3193 ; n3193_not
g30238 not n8620 ; n8620_not
g30239 not n4156 ; n4156_not
g30240 not n4525 ; n4525_not
g30241 not n2446 ; n2446_not
g30242 not n2275 ; n2275_not
g30243 not n5308 ; n5308_not
g30244 not n2239 ; n2239_not
g30245 not n5902 ; n5902_not
g30246 not n1933 ; n1933_not
g30247 not n5047 ; n5047_not
g30248 not n2653 ; n2653_not
g30249 not n1924 ; n1924_not
g30250 not n8611 ; n8611_not
g30251 not n5470 ; n5470_not
g30252 not n2455 ; n2455_not
g30253 not n1366 ; n1366_not
g30254 not n9160 ; n9160_not
g30255 not n5218 ; n5218_not
g30256 not n8431 ; n8431_not
g30257 not n4129 ; n4129_not
g30258 not n1357 ; n1357_not
g30259 not n7171 ; n7171_not
g30260 not n3364 ; n3364_not
g30261 not n4039 ; n4039_not
g30262 not n2266 ; n2266_not
g30263 not n2464 ; n2464_not
g30264 not n4507 ; n4507_not
g30265 not n5830 ; n5830_not
g30266 not n7162 ; n7162_not
g30267 not n3481 ; n3481_not
g30268 not n3175 ; n3175_not
g30269 not n4192 ; n4192_not
g30270 not n1294 ; n1294_not
g30271 not n7153 ; n7153_not
g30272 not n7036 ; n7036_not
g30273 not n5821 ; n5821_not
g30274 not n2851 ; n2851_not
g30275 not n3562 ; n3562_not
g30276 not n2635 ; n2635_not
g30277 not n9151 ; n9151_not
g30278 not n1267 ; n1267_not
g30279 not n4264 ; n4264_not
g30280 not n1942 ; n1942_not
g30281 not n5434 ; n5434_not
g30282 not n5227 ; n5227_not
g30283 not n4165 ; n4165_not
g30284 not n5029 ; n5029_not
g30285 not n8170 ; n8170_not
g30286 not n4174 ; n4174_not
g30287 not n1159 ; n1159_not
g30288 not n2626 ; n2626_not
g30289 not n3184 ; n3184_not
g30290 not n3436 ; n3436_not
g30291 not n6028 ; n6028_not
g30292 not n3508 ; n3508_not
g30293 not n4705 ; n4705_not
g30294 not n4480 ; n4480_not
g30295 not n4903 ; n4903_not
g30296 not n1744 ; n1744_not
g30297 not n5146 ; n5146_not
g30298 not n3760 ; n3760_not
g30299 not n1645 ; n1645_not
g30300 not n8305 ; n8305_not
g30301 not n6703 ; n6703_not
g30302 not n6802 ; n6802_not
g30303 not n9313 ; n9313_not
g30304 not n7513 ; n7513_not
g30305 not n4921 ; n4921_not
g30306 not n2392 ; n2392_not
g30307 not n8080 ; n8080_not
g30308 not n7081 ; n7081_not
g30309 not n2770 ; n2770_not
g30310 not n6640 ; n6640_not
g30311 not n6406 ; n6406_not
g30312 not n8440 ; n8440_not
g30313 not n5740 ; n5740_not
g30314 not n8062 ; n8062_not
g30315 not n7072 ; n7072_not
g30316 not n4723 ; n4723_not
g30317 not n1654 ; n1654_not
g30318 not n5506 ; n5506_not
g30319 not n3742 ; n3742_not
g30320 not n3634 ; n3634_not
g30321 not n9421 ; n9421_not
g30322 not n3058 ; n3058_not
g30323 not n2149 ; n2149_not
g30324 not n3391 ; n3391_not
g30325 not n7531 ; n7531_not
g30326 not n2545 ; n2545_not
g30327 not n4714 ; n4714_not
g30328 not n6523 ; n6523_not
g30329 not n6361 ; n6361_not
g30330 not n3373 ; n3373_not
g30331 not n7450 ; n7450_not
g30332 not n1636 ; n1636_not
g30333 not n5524 ; n5524_not
g30334 not n5155 ; n5155_not
g30335 not n2761 ; n2761_not
g30336 not n8350 ; n8350_not
g30337 not n4813 ; n4813_not
g30338 not n3805 ; n3805_not
g30339 not n6370 ; n6370_not
g30340 not n4660 ; n4660_not
g30341 not n6235 ; n6235_not
g30342 not n7090 ; n7090_not
g30343 not n1825 ; n1825_not
g30344 not n6712 ; n6712_not
g30345 not n4930 ; n4930_not
g30346 not n7504 ; n7504_not
g30347 not n3382 ; n3382_not
g30348 not n4390 ; n4390_not
g30349 not n1753 ; n1753_not
g30350 not n9304 ; n9304_not
g30351 not n1618 ; n1618_not
g30352 not n6721 ; n6721_not
g30353 not n2527 ; n2527_not
g30354 not n6730 ; n6730_not
g30355 not n6253 ; n6253_not
g30356 not n7423 ; n7423_not
g30357 not n9052 ; n9052_not
g30358 not n2536 ; n2536_not
g30359 not n1672 ; n1672_not
g30360 not n6604 ; n6604_not
g30361 not n7630 ; n7630_not
g30362 not n4417 ; n4417_not
g30363 not n7306 ; n7306_not
g30364 not n7621 ; n7621_not
g30365 not n8323 ; n8323_not
g30366 not n1681 ; n1681_not
g30367 not n2365 ; n2365_not
g30368 not n2167 ; n2167_not
g30369 not n6532 ; n6532_not
g30370 not n1708 ; n1708_not
g30371 not n4912 ; n4912_not
g30372 not n5335 ; n5335_not
g30373 not n5515 ; n5515_not
g30374 not n6622 ; n6622_not
g30375 not n3652 ; n3652_not
g30376 not n6244 ; n6244_not
g30377 not n6550 ; n6550_not
g30378 not n6181 ; n6181_not
g30379 not n4426 ; n4426_not
g30380 not n5119 ; n5119_not
g30381 not n3661 ; n3661_not
g30382 not n7702 ; n7702_not
g30383 not n7711 ; n7711_not
g30384 not n7720 ; n7720_not
g30385 not n3670 ; n3670_not
g30386 not n7342 ; n7342_not
g30387 not n8053 ; n8053_not
g30388 not n9403 ; n9403_not
g30389 not n3715 ; n3715_not
g30390 not n4750 ; n4750_not
g30391 not n4408 ; n4408_not
g30392 not n9412 ; n9412_not
g30393 not n9331 ; n9331_not
g30394 not n7261 ; n7261_not
g30395 not n1663 ; n1663_not
g30396 not n8314 ; n8314_not
g30397 not n4804 ; n4804_not
g30398 not n3724 ; n3724_not
g30399 not n4741 ; n4741_not
g30400 not n2176 ; n2176_not
g30401 not n1807 ; n1807_not
g30402 not n3733 ; n3733_not
g30403 not n6073 ; n6073_not
g30404 not n7603 ; n7603_not
g30405 not n6631 ; n6631_not
g30406 not n3418 ; n3418_not
g30407 not n6136 ; n6136_not
g30408 not n3643 ; n3643_not
g30409 not n9250 ; n9250_not
g30410 not n3706 ; n3706_not
g30411 not n5137 ; n5137_not
g30412 not n5128 ; n5128_not
g30413 not n5731 ; n5731_not
g30414 not n1546 ; n1546_not
g30415 not n9511 ; n9511_not
g30416 not n3904 ; n3904_not
g30417 not n2734 ; n2734_not
g30418 not n3607 ; n3607_not
g30419 not n4336 ; n4336_not
g30420 not n2329 ; n2329_not
g30421 not n1834 ; n1834_not
g30422 not n1852 ; n1852_not
g30423 not n2680 ; n2680_not
g30424 not n3463 ; n3463_not
g30425 not n2338 ; n2338_not
g30426 not n9232 ; n9232_not
g30427 not n8512 ; n8512_not
g30428 not n4732 ; n4732_not
g30429 not n2860 ; n2860_not
g30430 not n3328 ; n3328_not
g30431 not n1690 ; n1690_not
g30432 not n7333 ; n7333_not
g30433 not n1843 ; n1843_not
g30434 not n1582 ; n1582_not
g30435 not n6262 ; n6262_not
g30436 not n4606 ; n4606_not
g30437 not n7324 ; n7324_not
g30438 not n8044 ; n8044_not
g30439 not n7108 ; n7108_not
g30440 not n3319 ; n3319_not
g30441 not n9502 ; n9502_not
g30442 not n5074 ; n5074_not
g30443 not n4516 ; n4516_not
g30444 not n1555 ; n1555_not
g30445 not n6190 ; n6190_not
g30446 not n5605 ; n5605_not
g30447 not n7270 ; n7270_not
g30448 not n2725 ; n2725_not
g30449 not n1870 ; n1870_not
g30450 not n5254 ; n5254_not
g30451 not n7009 ; n7009_not
g30452 not n6343 ; n6343_not
g30453 not n3085 ; n3085_not
g30454 not n1474 ; n1474_not
g30455 not n9043 ; n9043_not
g30456 not n2716 ; n2716_not
g30457 not n4570 ; n4570_not
g30458 not n1735 ; n1735_not
g30459 not n3922 ; n3922_not
g30460 not n3913 ; n3913_not
g30461 not n6226 ; n6226_not
g30462 not n6019 ; n6019_not
g30463 not n6172 ; n6172_not
g30464 not n8152 ; n8152_not
g30465 not n6271 ; n6271_not
g30466 not n6910 ; n6910_not
g30467 not n4354 ; n4354_not
g30468 not n6280 ; n6280_not
g30469 not n3940 ; n3940_not
g30470 not n4444 ; n4444_not
g30471 not n3355 ; n3355_not
g30472 not n4435 ; n4435_not
g30473 not n5083 ; n5083_not
g30474 not n4642 ; n4642_not
g30475 not n6082 ; n6082_not
g30476 not n3517 ; n3517_not
g30477 not n7414 ; n7414_not
g30478 not n3841 ; n3841_not
g30479 not n4372 ; n4372_not
g30480 not n1591 ; n1591_not
g30481 not n3850 ; n3850_not
g30482 not n8503 ; n8503_not
g30483 not n6820 ; n6820_not
g30484 not n4633 ; n4633_not
g30485 not n5353 ; n5353_not
g30486 not n1609 ; n1609_not
g30487 not n3814 ; n3814_not
g30488 not n3067 ; n3067_not
g30489 not n3625 ; n3625_not
g30490 not n5380 ; n5380_not
g30491 not n9430 ; n9430_not
g30492 not n4651 ; n4651_not
g30493 not n7432 ; n7432_not
g30494 not n6352 ; n6352_not
g30495 not n6811 ; n6811_not
g30496 not n3832 ; n3832_not
g30497 not n6055 ; n6055_not
g30498 not n6046 ; n6046_not
g30499 not n7360 ; n7360_not
g30500 not n3337 ; n3337_not
g30501 not n7351 ; n7351_not
g30502 not n2914 ; n2914_not
g30503 not n5263 ; n5263_not
g30504 not n1771 ; n1771_not
g30505 not n2554 ; n2554_not
g30506 not n4624 ; n4624_not
g30507 not n8413 ; n8413_not
g30508 not n3616 ; n3616_not
g30509 not n3076 ; n3076_not
g30510 not n5038 ; n5038_not
g30511 not n2743 ; n2743_not
g30512 not n3346 ; n3346_not
g30513 not n4615 ; n4615_not
g30514 not n5164 ; n5164_not
g30515 not n2518 ; n2518_not
g30516 not n7405 ; n7405_not
g30517 not n5390 ; n5390_not
g30518 not n5255 ; n5255_not
g30519 not n5264 ; n5264_not
g30520 not n6425 ; n6425_not
g30521 not n5714 ; n5714_not
g30522 not n5543 ; n5543_not
g30523 not n5534 ; n5534_not
g30524 not n6443 ; n6443_not
g30525 not n5372 ; n5372_not
g30526 not n5345 ; n5345_not
g30527 not n4454 ; n4454_not
g30528 not n4472 ; n4472_not
g30529 not n6803 ; n6803_not
g30530 not n5750 ; n5750_not
g30531 not n6065 ; n6065_not
g30532 not n4238 ; n4238_not
g30533 not n4436 ; n4436_not
g30534 not n6128 ; n6128_not
g30535 not n5282 ; n5282_not
g30536 not n6173 ; n6173_not
g30537 not n6191 ; n6191_not
g30538 not n6182 ; n6182_not
g30539 not n7073 ; n7073_not
g30540 not n7055 ; n7055_not
g30541 not n4445 ; n4445_not
g30542 not n5057 ; n5057_not
g30543 not n4427 ; n4427_not
g30544 not n4733 ; n4733_not
g30545 not n5246 ; n5246_not
g30546 not n4463 ; n4463_not
g30547 not n6137 ; n6137_not
g30548 not n6434 ; n6434_not
g30549 not n5732 ; n5732_not
g30550 not n6290 ; n6290_not
g30551 not n6821 ; n6821_not
g30552 not n6083 ; n6083_not
g30553 not n4643 ; n4643_not
g30554 not n6254 ; n6254_not
g30555 not n4634 ; n4634_not
g30556 not n6812 ; n6812_not
g30557 not n5840 ; n5840_not
g30558 not n5525 ; n5525_not
g30559 not n6362 ; n6362_not
g30560 not n4652 ; n4652_not
g30561 not n4814 ; n4814_not
g30562 not n4940 ; n4940_not
g30563 not n5156 ; n5156_not
g30564 not n6371 ; n6371_not
g30565 not n4661 ; n4661_not
g30566 not n6731 ; n6731_not
g30567 not n6740 ; n6740_not
g30568 not n6722 ; n6722_not
g30569 not n4706 ; n4706_not
g30570 not n4580 ; n4580_not
g30571 not n6605 ; n6605_not
g30572 not n5606 ; n5606_not
g30573 not n6911 ; n6911_not
g30574 not n5552 ; n5552_not
g30575 not n5417 ; n5417_not
g30576 not n6272 ; n6272_not
g30577 not n6614 ; n6614_not
g30578 not n5480 ; n5480_not
g30579 not n6227 ; n6227_not
g30580 not n6092 ; n6092_not
g30581 not n5903 ; n5903_not
g30582 not n6047 ; n6047_not
g30583 not n5075 ; n5075_not
g30584 not n4616 ; n4616_not
g30585 not n6344 ; n6344_not
g30586 not n6056 ; n6056_not
g30587 not n4625 ; n4625_not
g30588 not n5165 ; n5165_not
g30589 not n4904 ; n4904_not
g30590 not n5516 ; n5516_not
g30591 not n6632 ; n6632_not
g30592 not n5570 ; n5570_not
g30593 not n5129 ; n5129_not
g30594 not n4913 ; n4913_not
g30595 not n6623 ; n6623_not
g30596 not n4760 ; n4760_not
g30597 not n4544 ; n4544_not
g30598 not n6335 ; n6335_not
g30599 not n6533 ; n6533_not
g30600 not n6038 ; n6038_not
g30601 not n5093 ; n5093_not
g30602 not n5336 ; n5336_not
g30603 not n4562 ; n4562_not
g30604 not n6326 ; n6326_not
g30605 not n6551 ; n6551_not
g30606 not n6713 ; n6713_not
g30607 not n4931 ; n4931_not
g30608 not n6380 ; n6380_not
g30609 not n6281 ; n6281_not
g30610 not n5138 ; n5138_not
g30611 not n5147 ; n5147_not
g30612 not n4715 ; n4715_not
g30613 not n6029 ; n6029_not
g30614 not n4724 ; n4724_not
g30615 not n6560 ; n6560_not
g30616 not n6407 ; n6407_not
g30617 not n6074 ; n6074_not
g30618 not n6650 ; n6650_not
g30619 not n6641 ; n6641_not
g30620 not n4805 ; n4805_not
g30621 not n4742 ; n4742_not
g30622 not n5741 ; n5741_not
g30623 not n6146 ; n6146_not
g30624 not n6155 ; n6155_not
g30625 not n5507 ; n5507_not
g30626 not n4517 ; n4517_not
g30627 not n6452 ; n6452_not
g30628 not n4526 ; n4526_not
g30629 not n6317 ; n6317_not
g30630 not n6245 ; n6245_not
g30631 not n5219 ; n5219_not
g30632 not n5660 ; n5660_not
g30633 not n5435 ; n5435_not
g30634 not n5318 ; n5318_not
g30635 not n6470 ; n6470_not
g30636 not n5048 ; n5048_not
g30637 not n5471 ; n5471_not
g30638 not n5408 ; n5408_not
g30639 not n5237 ; n5237_not
g30640 not n4481 ; n4481_not
g30641 not n7046 ; n7046_not
g30642 not n4490 ; n4490_not
g30643 not n5039 ; n5039_not
g30644 not n5291 ; n5291_not
g30645 not n6164 ; n6164_not
g30646 not n7037 ; n7037_not
g30647 not n5426 ; n5426_not
g30648 not n6119 ; n6119_not
g30649 not n5804 ; n5804_not
g30650 not n6461 ; n6461_not
g30651 not n5309 ; n5309_not
g30652 not n5813 ; n5813_not
g30653 not n5831 ; n5831_not
g30654 not n6308 ; n6308_not
g30655 not n5822 ; n5822_not
g30656 not n5705 ; n5705_not
g30657 not n5624 ; n5624_not
g30658 not n5462 ; n5462_not
g30659 not n5615 ; n5615_not
g30660 not n4823 ; n4823_not
g30661 not n4553 ; n4553_not
g30662 not n5183 ; n5183_not
g30663 not n7019 ; n7019_not
g30664 not n5327 ; n5327_not
g30665 not n6524 ; n6524_not
g30666 not n4571 ; n4571_not
g30667 not n5354 ; n5354_not
g30668 not n5066 ; n5066_not
g30669 not n5273 ; n5273_not
g30670 not n5651 ; n5651_not
g30671 not n7028 ; n7028_not
g30672 not n4841 ; n4841_not
g30673 not n5453 ; n5453_not
g30674 not n5912 ; n5912_not
g30675 not n5642 ; n5642_not
g30676 not n6506 ; n6506_not
g30677 not n5921 ; n5921_not
g30678 not n6209 ; n6209_not
g30679 not n5930 ; n5930_not
g30680 not n5633 ; n5633_not
g30681 not n5192 ; n5192_not
g30682 not n6416 ; n6416_not
g30683 not n6218 ; n6218_not
g30684 not n8243 ; n8243_not
g30685 not n2942 ; n2942_not
g30686 not n8252 ; n8252_not
g30687 not n2933 ; n2933_not
g30688 not n2744 ; n2744_not
g30689 not n2924 ; n2924_not
g30690 not n8261 ; n8261_not
g30691 not n8270 ; n8270_not
g30692 not n2915 ; n2915_not
g30693 not n2861 ; n2861_not
g30694 not n2906 ; n2906_not
g30695 not n8306 ; n8306_not
g30696 not n8324 ; n8324_not
g30697 not n2870 ; n2870_not
g30698 not n8342 ; n8342_not
g30699 not n8351 ; n8351_not
g30700 not n8360 ; n8360_not
g30701 not n8081 ; n8081_not
g30702 not n2852 ; n2852_not
g30703 not n3158 ; n3158_not
g30704 not n3149 ; n3149_not
g30705 not n3095 ; n3095_not
g30706 not n8144 ; n8144_not
g30707 not n3086 ; n3086_not
g30708 not n3077 ; n3077_not
g30709 not n3068 ; n3068_not
g30710 not n3059 ; n3059_not
g30711 not n8153 ; n8153_not
g30712 not n8171 ; n8171_not
g30713 not n8207 ; n8207_not
g30714 not n2654 ; n2654_not
g30715 not n8216 ; n8216_not
g30716 not n8018 ; n8018_not
g30717 not n8225 ; n8225_not
g30718 not n2951 ; n2951_not
g30719 not n2960 ; n2960_not
g30720 not n8234 ; n8234_not
g30721 not n2735 ; n2735_not
g30722 not n8513 ; n8513_not
g30723 not n2717 ; n2717_not
g30724 not n2726 ; n2726_not
g30725 not n2708 ; n2708_not
g30726 not n8522 ; n8522_not
g30727 not n2690 ; n2690_not
g30728 not n8531 ; n8531_not
g30729 not n2681 ; n2681_not
g30730 not n2555 ; n2555_not
g30731 not n2663 ; n2663_not
g30732 not n8603 ; n8603_not
g30733 not n8612 ; n8612_not
g30734 not n2645 ; n2645_not
g30735 not n2492 ; n2492_not
g30736 not n2636 ; n2636_not
g30737 not n8621 ; n8621_not
g30738 not n2627 ; n2627_not
g30739 not n2618 ; n2618_not
g30740 not n2843 ; n2843_not
g30741 not n2834 ; n2834_not
g30742 not n2816 ; n2816_not
g30743 not n2807 ; n2807_not
g30744 not n2483 ; n2483_not
g30745 not n8414 ; n8414_not
g30746 not n8423 ; n8423_not
g30747 not n2780 ; n2780_not
g30748 not n8441 ; n8441_not
g30749 not n2771 ; n2771_not
g30750 not n8450 ; n8450_not
g30751 not n2762 ; n2762_not
g30752 not n8315 ; n8315_not
g30753 not n2753 ; n2753_not
g30754 not n8504 ; n8504_not
g30755 not n7460 ; n7460_not
g30756 not n7802 ; n7802_not
g30757 not n7811 ; n7811_not
g30758 not n3590 ; n3590_not
g30759 not n7820 ; n7820_not
g30760 not n3581 ; n3581_not
g30761 not n7910 ; n7910_not
g30762 not n3572 ; n3572_not
g30763 not n7721 ; n7721_not
g30764 not n3563 ; n3563_not
g30765 not n3554 ; n3554_not
g30766 not n3545 ; n3545_not
g30767 not n3536 ; n3536_not
g30768 not n3527 ; n3527_not
g30769 not n3518 ; n3518_not
g30770 not n3509 ; n3509_not
g30771 not n3491 ; n3491_not
g30772 not n3734 ; n3734_not
g30773 not n3725 ; n3725_not
g30774 not n3716 ; n3716_not
g30775 not n7604 ; n7604_not
g30776 not n3482 ; n3482_not
g30777 not n7622 ; n7622_not
g30778 not n3680 ; n3680_not
g30779 not n3473 ; n3473_not
g30780 not n7640 ; n7640_not
g30781 not n3671 ; n3671_not
g30782 not n7712 ; n7712_not
g30783 not n3653 ; n3653_not
g30784 not n3617 ; n3617_not
g30785 not n7730 ; n7730_not
g30786 not n3644 ; n3644_not
g30787 not n3635 ; n3635_not
g30788 not n3437 ; n3437_not
g30789 not n3626 ; n3626_not
g30790 not n3455 ; n3455_not
g30791 not n3338 ; n3338_not
g30792 not n8108 ; n8108_not
g30793 not n3293 ; n3293_not
g30794 not n8117 ; n8117_not
g30795 not n3275 ; n3275_not
g30796 not n3284 ; n3284_not
g30797 not n3266 ; n3266_not
g30798 not n3257 ; n3257_not
g30799 not n3248 ; n3248_not
g30800 not n3239 ; n3239_not
g30801 not n3176 ; n3176_not
g30802 not n8126 ; n8126_not
g30803 not n3194 ; n3194_not
g30804 not n3185 ; n3185_not
g30805 not n8054 ; n8054_not
g30806 not n3167 ; n3167_not
g30807 not n8135 ; n8135_not
g30808 not n8027 ; n8027_not
g30809 not n3464 ; n3464_not
g30810 not n8045 ; n8045_not
g30811 not n3446 ; n3446_not
g30812 not n3428 ; n3428_not
g30813 not n3419 ; n3419_not
g30814 not n3356 ; n3356_not
g30815 not n8063 ; n8063_not
g30816 not n3392 ; n3392_not
g30817 not n3374 ; n3374_not
g30818 not n3365 ; n3365_not
g30819 not n3347 ; n3347_not
g30820 not n9071 ; n9071_not
g30821 not n1718 ; n1718_not
g30822 not n1709 ; n1709_not
g30823 not n9350 ; n9350_not
g30824 not n1691 ; n1691_not
g30825 not n9305 ; n9305_not
g30826 not n1682 ; n1682_not
g30827 not n9404 ; n9404_not
g30828 not n1673 ; n1673_not
g30829 not n1664 ; n1664_not
g30830 not n9422 ; n9422_not
g30831 not n1646 ; n1646_not
g30832 not n1637 ; n1637_not
g30833 not n1628 ; n1628_not
g30834 not n1619 ; n1619_not
g30835 not n9431 ; n9431_not
g30836 not n9440 ; n9440_not
g30837 not n1592 ; n1592_not
g30838 not n9152 ; n9152_not
g30839 not n9224 ; n9224_not
g30840 not n1862 ; n1862_not
g30841 not n1853 ; n1853_not
g30842 not n9233 ; n9233_not
g30843 not n1844 ; n1844_not
g30844 not n1835 ; n1835_not
g30845 not n9251 ; n9251_not
g30846 not n9260 ; n9260_not
g30847 not n1745 ; n1745_not
g30848 not n1817 ; n1817_not
g30849 not n1808 ; n1808_not
g30850 not n1772 ; n1772_not
g30851 not n9314 ; n9314_not
g30852 not n1754 ; n1754_not
g30853 not n9332 ; n9332_not
g30854 not n1736 ; n1736_not
g30855 not n9701 ; n9701_not
g30856 not n1358 ; n1358_not
g30857 not n1268 ; n1268_not
g30858 not n9800 ; n9800_not
g30859 not n1295 ; n1295_not
g30860 not n1277 ; n1277_not
g30861 not n1259 ; n1259_not
g30862 not n1196 ; n1196_not
g30863 not n1187 ; n1187_not
g30864 not n1178 ; n1178_not
g30865 not n1169 ; n1169_not
g30866 not n7703 ; n7703_not
g30867 not n1088 ; n1088_not
g30868 not n1097 ; n1097_not
g30869 not n1079 ; n1079_not
g30870 not n6515 ; n6515_not
g30871 not n4922 ; n4922_not
g30872 not n3383 ; n3383_not
g30873 not n9503 ; n9503_not
g30874 not n1583 ; n1583_not
g30875 not n9512 ; n9512_not
g30876 not n1574 ; n1574_not
g30877 not n1565 ; n1565_not
g30878 not n9530 ; n9530_not
g30879 not n1556 ; n1556_not
g30880 not n1547 ; n1547_not
g30881 not n1538 ; n1538_not
g30882 not n1493 ; n1493_not
g30883 not n1484 ; n1484_not
g30884 not n1475 ; n1475_not
g30885 not n9611 ; n9611_not
g30886 not n1448 ; n1448_not
g30887 not n1457 ; n1457_not
g30888 not n1439 ; n1439_not
g30889 not n1385 ; n1385_not
g30890 not n1376 ; n1376_not
g30891 not n2465 ; n2465_not
g30892 not n2456 ; n2456_not
g30893 not n8900 ; n8900_not
g30894 not n2447 ; n2447_not
g30895 not n2429 ; n2429_not
g30896 not n2339 ; n2339_not
g30897 not n2393 ; n2393_not
g30898 not n2384 ; n2384_not
g30899 not n2375 ; n2375_not
g30900 not n2366 ; n2366_not
g30901 not n9017 ; n9017_not
g30902 not n2357 ; n2357_not
g30903 not n2348 ; n2348_not
g30904 not n2249 ; n2249_not
g30905 not n2294 ; n2294_not
g30906 not n2609 ; n2609_not
g30907 not n8630 ; n8630_not
g30908 not n2582 ; n2582_not
g30909 not n2591 ; n2591_not
g30910 not n8702 ; n8702_not
g30911 not n2573 ; n2573_not
g30912 not n2564 ; n2564_not
g30913 not n8720 ; n8720_not
g30914 not n2546 ; n2546_not
g30915 not n2537 ; n2537_not
g30916 not n2528 ; n2528_not
g30917 not n2519 ; n2519_not
g30918 not n8711 ; n8711_not
g30919 not n8405 ; n8405_not
g30920 not n8801 ; n8801_not
g30921 not n2474 ; n2474_not
g30922 not n9116 ; n9116_not
g30923 not n9044 ; n9044_not
g30924 not n9125 ; n9125_not
g30925 not n1970 ; n1970_not
g30926 not n1961 ; n1961_not
g30927 not n1952 ; n1952_not
g30928 not n9143 ; n9143_not
g30929 not n1943 ; n1943_not
g30930 not n9161 ; n9161_not
g30931 not n1934 ; n1934_not
g30932 not n1925 ; n1925_not
g30933 not n1916 ; n1916_not
g30934 not n9008 ; n9008_not
g30935 not n1880 ; n1880_not
g30936 not n9215 ; n9215_not
g30937 not n1871 ; n1871_not
g30938 not n2285 ; n2285_not
g30939 not n9035 ; n9035_not
g30940 not n2276 ; n2276_not
g30941 not n2267 ; n2267_not
g30942 not n2258 ; n2258_not
g30943 not n2195 ; n2195_not
g30944 not n2177 ; n2177_not
g30945 not n2168 ; n2168_not
g30946 not n2159 ; n2159_not
g30947 not n9053 ; n9053_not
g30948 not n2087 ; n2087_not
g30949 not n2078 ; n2078_not
g30950 not n2069 ; n2069_not
g30951 not n9107 ; n9107_not
g30952 not n7343 ; n7343_not
g30953 not n7325 ; n7325_not
g30954 not n3905 ; n3905_not
g30955 not n3914 ; n3914_not
g30956 not n3923 ; n3923_not
g30957 not n7307 ; n7307_not
g30958 not n3932 ; n3932_not
g30959 not n3941 ; n3941_not
g30960 not n7280 ; n7280_not
g30961 not n7271 ; n7271_not
g30962 not n3950 ; n3950_not
g30963 not n7262 ; n7262_not
g30964 not n7253 ; n7253_not
g30965 not n7244 ; n7244_not
g30966 not n3824 ; n3824_not
g30967 not n7235 ; n7235_not
g30968 not n7217 ; n7217_not
g30969 not n4049 ; n4049_not
g30970 not n4067 ; n4067_not
g30971 not n4094 ; n4094_not
g30972 not n7523 ; n7523_not
g30973 not n3761 ; n3761_not
g30974 not n7514 ; n7514_not
g30975 not n7505 ; n7505_not
g30976 not n7451 ; n7451_not
g30977 not n3806 ; n3806_not
g30978 not n7442 ; n7442_not
g30979 not n3815 ; n3815_not
g30980 not n7433 ; n7433_not
g30981 not n3833 ; n3833_not
g30982 not n7424 ; n7424_not
g30983 not n7415 ; n7415_not
g30984 not n3851 ; n3851_not
g30985 not n7406 ; n7406_not
g30986 not n7370 ; n7370_not
g30987 not n7352 ; n7352_not
g30988 not n4283 ; n4283_not
g30989 not n4292 ; n4292_not
g30990 not n7118 ; n7118_not
g30991 not n4328 ; n4328_not
g30992 not n4319 ; n4319_not
g30993 not n4337 ; n4337_not
g30994 not n4346 ; n4346_not
g30995 not n4355 ; n4355_not
g30996 not n7109 ; n7109_not
g30997 not n4364 ; n4364_not
g30998 not n4373 ; n4373_not
g30999 not n7091 ; n7091_not
g31000 not n7082 ; n7082_not
g31001 not n4391 ; n4391_not
g31002 not n4409 ; n4409_not
g31003 not n4418 ; n4418_not
g31004 not n7190 ; n7190_not
g31005 not n7181 ; n7181_not
g31006 not n4139 ; n4139_not
g31007 not n4148 ; n4148_not
g31008 not n4157 ; n4157_not
g31009 not n4166 ; n4166_not
g31010 not n4175 ; n4175_not
g31011 not n7172 ; n7172_not
g31012 not n4184 ; n4184_not
g31013 not n7163 ; n7163_not
g31014 not n7154 ; n7154_not
g31015 not n4229 ; n4229_not
g31016 not n4247 ; n4247_not
g31017 not n7145 ; n7145_not
g31018 not n4256 ; n4256_not
g31019 not n4265 ; n4265_not
g31020 not n7136 ; n7136_not
g31021 not n4274 ; n4274_not
g31022 not n7127 ; n7127_not
g31023 not n3743 ; n3743_not
g31024 not n7550 ; n7550_not
g31025 not n7532 ; n7532_not
g31026 not n3752 ; n3752_not
g31027 not n4059 ; n4059_not
g31028 not n2268 ; n2268_not
g31029 not n7371 ; n7371_not
g31030 not n6129 ; n6129_not
g31031 not n2169 ; n2169_not
g31032 not n2259 ; n2259_not
g31033 not n4068 ; n4068_not
g31034 not n4077 ; n4077_not
g31035 not n7137 ; n7137_not
g31036 not n4086 ; n4086_not
g31037 not n2196 ; n2196_not
g31038 not n5373 ; n5373_not
g31039 not n9054 ; n9054_not
g31040 not n2187 ; n2187_not
g31041 not n2178 ; n2178_not
g31042 not n7191 ; n7191_not
g31043 not n6138 ; n6138_not
g31044 not n7029 ; n7029_not
g31045 not n1980 ; n1980_not
g31046 not n1971 ; n1971_not
g31047 not n7236 ; n7236_not
g31048 not n2376 ; n2376_not
g31049 not n2367 ; n2367_not
g31050 not n4554 ; n4554_not
g31051 not n2358 ; n2358_not
g31052 not n9018 ; n9018_not
g31053 not n7227 ; n7227_not
g31054 not n2349 ; n2349_not
g31055 not n5346 ; n5346_not
g31056 not n7218 ; n7218_not
g31057 not n6156 ; n6156_not
g31058 not n7704 ; n7704_not
g31059 not n9027 ; n9027_not
g31060 not n2295 ; n2295_not
g31061 not n2286 ; n2286_not
g31062 not n7209 ; n7209_not
g31063 not n5355 ; n5355_not
g31064 not n6147 ; n6147_not
g31065 not n9036 ; n9036_not
g31066 not n2277 ; n2277_not
g31067 not n3663 ; n3663_not
g31068 not n5364 ; n5364_not
g31069 not n9135 ; n9135_not
g31070 not n1962 ; n1962_not
g31071 not n5427 ; n5427_not
g31072 not n4167 ; n4167_not
g31073 not n4518 ; n4518_not
g31074 not n7173 ; n7173_not
g31075 not n9144 ; n9144_not
g31076 not n1872 ; n1872_not
g31077 not n1944 ; n1944_not
g31078 not n6660 ; n6660_not
g31079 not n4176 ; n4176_not
g31080 not n5436 ; n5436_not
g31081 not n1935 ; n1935_not
g31082 not n6606 ; n6606_not
g31083 not n1926 ; n1926_not
g31084 not n9162 ; n9162_not
g31085 not n9153 ; n9153_not
g31086 not n9171 ; n9171_not
g31087 not n5445 ; n5445_not
g31088 not n9009 ; n9009_not
g31089 not n9180 ; n9180_not
g31090 not n5454 ; n5454_not
g31091 not n9207 ; n9207_not
g31092 not n9063 ; n9063_not
g31093 not n2097 ; n2097_not
g31094 not n2088 ; n2088_not
g31095 not n7542 ; n7542_not
g31096 not n2079 ; n2079_not
g31097 not n4095 ; n4095_not
g31098 not n3672 ; n3672_not
g31099 not n9072 ; n9072_not
g31100 not n9081 ; n9081_not
g31101 not n9090 ; n9090_not
g31102 not n5409 ; n5409_not
g31103 not n4149 ; n4149_not
g31104 not n9108 ; n9108_not
g31105 not n9117 ; n9117_not
g31106 not n5247 ; n5247_not
g31107 not n9045 ; n9045_not
g31108 not n4158 ; n4158_not
g31109 not n5418 ; n5418_not
g31110 not n9126 ; n9126_not
g31111 not n1827 ; n1827_not
g31112 not n2628 ; n2628_not
g31113 not n2637 ; n2637_not
g31114 not n5157 ; n5157_not
g31115 not n6921 ; n6921_not
g31116 not n7290 ; n7290_not
g31117 not n2619 ; n2619_not
g31118 not n6930 ; n6930_not
g31119 not n8622 ; n8622_not
g31120 not n4527 ; n4527_not
g31121 not n8613 ; n8613_not
g31122 not n8631 ; n8631_not
g31123 not n5238 ; n5238_not
g31124 not n2592 ; n2592_not
g31125 not n4581 ; n4581_not
g31126 not n8640 ; n8640_not
g31127 not n2583 ; n2583_not
g31128 not n8703 ; n8703_not
g31129 not n2574 ; n2574_not
g31130 not n8361 ; n8361_not
g31131 not n7281 ; n7281_not
g31132 not n5256 ; n5256_not
g31133 not n2565 ; n2565_not
g31134 not n5184 ; n5184_not
g31135 not n2709 ; n2709_not
g31136 not n3924 ; n3924_not
g31137 not n8523 ; n8523_not
g31138 not n2691 ; n2691_not
g31139 not n7308 ; n7308_not
g31140 not n8532 ; n8532_not
g31141 not n6903 ; n6903_not
g31142 not n2538 ; n2538_not
g31143 not n7533 ; n7533_not
g31144 not n2529 ; n2529_not
g31145 not n8550 ; n8550_not
g31146 not n8253 ; n8253_not
g31147 not n2664 ; n2664_not
g31148 not n3654 ; n3654_not
g31149 not n3933 ; n3933_not
g31150 not n6543 ; n6543_not
g31151 not n8604 ; n8604_not
g31152 not n2646 ; n2646_not
g31153 not n6912 ; n6912_not
g31154 not n8802 ; n8802_not
g31155 not n8811 ; n8811_not
g31156 not n2484 ; n2484_not
g31157 not n8820 ; n8820_not
g31158 not n3960 ; n3960_not
g31159 not n5274 ; n5274_not
g31160 not n2475 ; n2475_not
g31161 not n6354 ; n6354_not
g31162 not n2466 ; n2466_not
g31163 not n4563 ; n4563_not
g31164 not n8901 ; n8901_not
g31165 not n2457 ; n2457_not
g31166 not n5319 ; n5319_not
g31167 not n7254 ; n7254_not
g31168 not n8910 ; n8910_not
g31169 not n2448 ; n2448_not
g31170 not n2439 ; n2439_not
g31171 not n5328 ; n5328_not
g31172 not n7245 ; n7245_not
g31173 not n6570 ; n6570_not
g31174 not n2385 ; n2385_not
g31175 not n4545 ; n4545_not
g31176 not n5067 ; n5067_not
g31177 not n8721 ; n8721_not
g31178 not n2556 ; n2556_not
g31179 not n6192 ; n6192_not
g31180 not n2547 ; n2547_not
g31181 not n7272 ; n7272_not
g31182 not n5049 ; n5049_not
g31183 not n8730 ; n8730_not
g31184 not n3825 ; n3825_not
g31185 not n5283 ; n5283_not
g31186 not n6174 ; n6174_not
g31187 not n3951 ; n3951_not
g31188 not n7713 ; n7713_not
g31189 not n8712 ; n8712_not
g31190 not n2493 ; n2493_not
g31191 not n5292 ; n5292_not
g31192 not n4572 ; n4572_not
g31193 not n6165 ; n6165_not
g31194 not n1494 ; n1494_not
g31195 not n5625 ; n5625_not
g31196 not n5940 ; n5940_not
g31197 not n4338 ; n4338_not
g31198 not n6633 ; n6633_not
g31199 not n4356 ; n4356_not
g31200 not n5931 ; n5931_not
g31201 not n1476 ; n1476_not
g31202 not n9612 ; n9612_not
g31203 not n5913 ; n5913_not
g31204 not n5922 ; n5922_not
g31205 not n5472 ; n5472_not
g31206 not n6642 ; n6642_not
g31207 not n9630 ; n9630_not
g31208 not n1458 ; n1458_not
g31209 not n5643 ; n5643_not
g31210 not n4365 ; n4365_not
g31211 not n1449 ; n1449_not
g31212 not n4743 ; n4743_not
g31213 not n1386 ; n1386_not
g31214 not n5652 ; n5652_not
g31215 not n4446 ; n4446_not
g31216 not n5904 ; n5904_not
g31217 not n4266 ; n4266_not
g31218 not n9450 ; n9450_not
g31219 not n9504 ; n9504_not
g31220 not n4329 ; n4329_not
g31221 not n9513 ; n9513_not
g31222 not n1575 ; n1575_not
g31223 not n7056 ; n7056_not
g31224 not n3735 ; n3735_not
g31225 not n9522 ; n9522_not
g31226 not n6561 ; n6561_not
g31227 not n1557 ; n1557_not
g31228 not n4455 ; n4455_not
g31229 not n5607 ; n5607_not
g31230 not n9531 ; n9531_not
g31231 not n1548 ; n1548_not
g31232 not n3717 ; n3717_not
g31233 not n1485 ; n1485_not
g31234 not n1539 ; n1539_not
g31235 not n4347 ; n4347_not
g31236 not n5616 ; n5616_not
g31237 not n5805 ; n5805_not
g31238 not n4392 ; n4392_not
g31239 not n9900 ; n9900_not
g31240 not n1197 ; n1197_not
g31241 not n4437 ; n4437_not
g31242 not n1179 ; n1179_not
g31243 not n1188 ; n1188_not
g31244 not n7074 ; n7074_not
g31245 not n5706 ; n5706_not
g31246 not n9342 ; n9342_not
g31247 not n4239 ; n4239_not
g31248 not n1098 ; n1098_not
g31249 not n5715 ; n5715_not
g31250 not n5526 ; n5526_not
g31251 not n5751 ; n5751_not
g31252 not n7551 ; n7551_not
g31253 not n1089 ; n1089_not
g31254 not n4428 ; n4428_not
g31255 not n4419 ; n4419_not
g31256 not n5733 ; n5733_not
g31257 not n1377 ; n1377_not
g31258 not n4374 ; n4374_not
g31259 not n1359 ; n1359_not
g31260 not n4383 ; n4383_not
g31261 not n5661 ; n5661_not
g31262 not n9702 ; n9702_not
g31263 not n5850 ; n5850_not
g31264 not n5841 ; n5841_not
g31265 not n9711 ; n9711_not
g31266 not n5742 ; n5742_not
g31267 not n7083 ; n7083_not
g31268 not n5832 ; n5832_not
g31269 not n1296 ; n1296_not
g31270 not n4608 ; n4608_not
g31271 not n9801 ; n9801_not
g31272 not n5823 ; n5823_not
g31273 not n9810 ; n9810_not
g31274 not n5814 ; n5814_not
g31275 not n1287 ; n1287_not
g31276 not n1278 ; n1278_not
g31277 not n1269 ; n1269_not
g31278 not n6615 ; n6615_not
g31279 not n1683 ; n1683_not
g31280 not n4248 ; n4248_not
g31281 not n9261 ; n9261_not
g31282 not n7146 ; n7146_not
g31283 not n7614 ; n7614_not
g31284 not n1746 ; n1746_not
g31285 not n9270 ; n9270_not
g31286 not n1809 ; n1809_not
g31287 not n6075 ; n6075_not
g31288 not n5508 ; n5508_not
g31289 not n5517 ; n5517_not
g31290 not n1791 ; n1791_not
g31291 not n9306 ; n9306_not
g31292 not n1782 ; n1782_not
g31293 not n1773 ; n1773_not
g31294 not n3690 ; n3690_not
g31295 not n4761 ; n4761_not
g31296 not n7164 ; n7164_not
g31297 not n1881 ; n1881_not
g31298 not n7623 ; n7623_not
g31299 not n9216 ; n9216_not
g31300 not n7155 ; n7155_not
g31301 not n9225 ; n9225_not
g31302 not n4194 ; n4194_not
g31303 not n1863 ; n1863_not
g31304 not n1854 ; n1854_not
g31305 not n9234 ; n9234_not
g31306 not n5481 ; n5481_not
g31307 not n6093 ; n6093_not
g31308 not n9243 ; n9243_not
g31309 not n1845 ; n1845_not
g31310 not n1836 ; n1836_not
g31311 not n6084 ; n6084_not
g31312 not n9252 ; n9252_not
g31313 not n1692 ; n1692_not
g31314 not n5562 ; n5562_not
g31315 not n6039 ; n6039_not
g31316 not n4473 ; n4473_not
g31317 not n9405 ; n9405_not
g31318 not n1665 ; n1665_not
g31319 not n5571 ; n5571_not
g31320 not n7128 ; n7128_not
g31321 not n6651 ; n6651_not
g31322 not n1593 ; n1593_not
g31323 not n1647 ; n1647_not
g31324 not n4293 ; n4293_not
g31325 not n1638 ; n1638_not
g31326 not n3708 ; n3708_not
g31327 not n7119 ; n7119_not
g31328 not n5580 ; n5580_not
g31329 not n9441 ; n9441_not
g31330 not n4464 ; n4464_not
g31331 not n3681 ; n3681_not
g31332 not n9315 ; n9315_not
g31333 not n1764 ; n1764_not
g31334 not n6066 ; n6066_not
g31335 not n9324 ; n9324_not
g31336 not n1755 ; n1755_not
g31337 not n7605 ; n7605_not
g31338 not n7047 ; n7047_not
g31339 not n5535 ; n5535_not
g31340 not n4275 ; n4275_not
g31341 not n9333 ; n9333_not
g31342 not n1737 ; n1737_not
g31343 not n5544 ; n5544_not
g31344 not n6057 ; n6057_not
g31345 not n4482 ; n4482_not
g31346 not n1719 ; n1719_not
g31347 not n4284 ; n4284_not
g31348 not n6624 ; n6624_not
g31349 not n9351 ; n9351_not
g31350 not n5553 ; n5553_not
g31351 not n9360 ; n9360_not
g31352 not n3447 ; n3447_not
g31353 not n8226 ; n8226_not
g31354 not n3780 ; n3780_not
g31355 not n3456 ; n3456_not
g31356 not n8046 ; n8046_not
g31357 not n6417 ; n6417_not
g31358 not n3636 ; n3636_not
g31359 not n2961 ; n2961_not
g31360 not n2952 ; n2952_not
g31361 not n8235 ; n8235_not
g31362 not n2763 ; n2763_not
g31363 not n7407 ; n7407_not
g31364 not n8244 ; n8244_not
g31365 not n5058 ; n5058_not
g31366 not n2943 ; n2943_not
g31367 not n4680 ; n4680_not
g31368 not n8064 ; n8064_not
g31369 not n8172 ; n8172_not
g31370 not n3393 ; n3393_not
g31371 not n3573 ; n3573_not
g31372 not n8190 ; n8190_not
g31373 not n3294 ; n3294_not
g31374 not n3834 ; n3834_not
g31375 not n8208 ; n8208_not
g31376 not n6813 ; n6813_not
g31377 not n3429 ; n3429_not
g31378 not n4644 ; n4644_not
g31379 not n2970 ; n2970_not
g31380 not n3438 ; n3438_not
g31381 not n4905 ; n4905_not
g31382 not n2916 ; n2916_not
g31383 not n6714 ; n6714_not
g31384 not n3483 ; n3483_not
g31385 not n3564 ; n3564_not
g31386 not n6822 ; n6822_not
g31387 not n8019 ; n8019_not
g31388 not n8280 ; n8280_not
g31389 not n2907 ; n2907_not
g31390 not n6255 ; n6255_not
g31391 not n6426 ; n6426_not
g31392 not n8307 ; n8307_not
g31393 not n7506 ; n7506_not
g31394 not n3519 ; n3519_not
g31395 not n8316 ; n8316_not
g31396 not n2880 ; n2880_not
g31397 not n3771 ; n3771_not
g31398 not n8325 ; n8325_not
g31399 not n5094 ; n5094_not
g31400 not n4635 ; n4635_not
g31401 not n7740 ; n7740_not
g31402 not n3852 ; n3852_not
g31403 not n2934 ; n2934_not
g31404 not n4806 ; n4806_not
g31405 not n8262 ; n8262_not
g31406 not n8037 ; n8037_not
g31407 not n6273 ; n6273_not
g31408 not n2925 ; n2925_not
g31409 not n3474 ; n3474_not
g31410 not n7911 ; n7911_not
g31411 not n8271 ; n8271_not
g31412 not n8028 ; n8028_not
g31413 not n5076 ; n5076_not
g31414 not n6741 ; n6741_not
g31415 not n4941 ; n4941_not
g31416 not n3258 ; n3258_not
g31417 not n3249 ; n3249_not
g31418 not n7452 ; n7452_not
g31419 not n3069 ; n3069_not
g31420 not n4662 ; n4662_not
g31421 not n8127 ; n8127_not
g31422 not n3195 ; n3195_not
g31423 not n3177 ; n3177_not
g31424 not n3366 ; n3366_not
g31425 not n4716 ; n4716_not
g31426 not n8055 ; n8055_not
g31427 not n3186 ; n3186_not
g31428 not n3618 ; n3618_not
g31429 not n6336 ; n6336_not
g31430 not n6345 ; n6345_not
g31431 not n6534 ; n6534_not
g31432 not n7425 ; n7425_not
g31433 not n6750 ; n6750_not
g31434 not n7461 ; n7461_not
g31435 not n3357 ; n3357_not
g31436 not n6246 ; n6246_not
g31437 not n3285 ; n3285_not
g31438 not n4671 ; n4671_not
g31439 not n3276 ; n3276_not
g31440 not n8118 ; n8118_not
g31441 not n3267 ; n3267_not
g31442 not n8109 ; n8109_not
g31443 not n6327 ; n6327_not
g31444 not n6363 ; n6363_not
g31445 not n4653 ; n4653_not
g31446 not n3087 ; n3087_not
g31447 not n7434 ; n7434_not
g31448 not n3627 ; n3627_not
g31449 not n6291 ; n6291_not
g31450 not n6381 ; n6381_not
g31451 not n8145 ; n8145_not
g31452 not n6390 ; n6390_not
g31453 not n6282 ; n6282_not
g31454 not n8082 ; n8082_not
g31455 not n6732 ; n6732_not
g31456 not n4923 ; n4923_not
g31457 not n8154 ; n8154_not
g31458 not n8073 ; n8073_not
g31459 not n2826 ; n2826_not
g31460 not n8163 ; n8163_not
g31461 not n6309 ; n6309_not
g31462 not n7812 ; n7812_not
g31463 not n7470 ; n7470_not
g31464 not n3807 ; n3807_not
g31465 not n4815 ; n4815_not
g31466 not n3168 ; n3168_not
g31467 not n4491 ; n4491_not
g31468 not n6372 ; n6372_not
g31469 not n3159 ; n3159_not
g31470 not n4932 ; n4932_not
g31471 not n6804 ; n6804_not
g31472 not n8136 ; n8136_not
g31473 not n7443 ; n7443_not
g31474 not n8091 ; n8091_not
g31475 not n3384 ; n3384_not
g31476 not n3096 ; n3096_not
g31477 not n6840 ; n6840_not
g31478 not n5139 ; n5139_not
g31479 not n4851 ; n4851_not
g31480 not n8433 ; n8433_not
g31481 not n7920 ; n7920_not
g31482 not n8442 ; n8442_not
g31483 not n5148 ; n5148_not
g31484 not n2772 ; n2772_not
g31485 not n7326 ; n7326_not
g31486 not n7731 ; n7731_not
g31487 not n4734 ; n4734_not
g31488 not n4842 ; n4842_not
g31489 not n7524 ; n7524_not
g31490 not n4617 ; n4617_not
g31491 not n8406 ; n8406_not
g31492 not n2808 ; n2808_not
g31493 not n7344 ; n7344_not
g31494 not n3645 ; n3645_not
g31495 not n8415 ; n8415_not
g31496 not n7515 ; n7515_not
g31497 not n7722 ; n7722_not
g31498 not n6471 ; n6471_not
g31499 not n2790 ; n2790_not
g31500 not n3753 ; n3753_not
g31501 not n2781 ; n2781_not
g31502 not n6480 ; n6480_not
g31503 not n3906 ; n3906_not
g31504 not n8505 ; n8505_not
g31505 not n2736 ; n2736_not
g31506 not n6516 ; n6516_not
g31507 not n4590 ; n4590_not
g31508 not n3915 ; n3915_not
g31509 not n2727 ; n2727_not
g31510 not n4824 ; n4824_not
g31511 not n5175 ; n5175_not
g31512 not n2718 ; n2718_not
g31513 not n8514 ; n8514_not
g31514 not n2682 ; n2682_not
g31515 not n7803 ; n7803_not
g31516 not n2655 ; n2655_not
g31517 not n8460 ; n8460_not
g31518 not n4950 ; n4950_not
g31519 not n3582 ; n3582_not
g31520 not n2754 ; n2754_not
g31521 not n7902 ; n7902_not
g31522 not n2745 ; n2745_not
g31523 not n7317 ; n7317_not
g31524 not n5166 ; n5166_not
g31525 not n7821 ; n7821_not
g31526 not n4707 ; n4707_not
g31527 not n6228 ; n6228_not
g31528 not n2844 ; n2844_not
g31529 not n8343 ; n8343_not
g31530 not n7380 ; n7380_not
g31531 not n3528 ; n3528_not
g31532 not n4860 ; n4860_not
g31533 not n6705 ; n6705_not
g31534 not n3537 ; n3537_not
g31535 not n2862 ; n2862_not
g31536 not n8352 ; n8352_not
g31537 not n6462 ; n6462_not
g31538 not n6444 ; n6444_not
g31539 not n3555 ; n3555_not
g31540 not n3762 ; n3762_not
g31541 not n3744 ; n3744_not
g31542 not n8370 ; n8370_not
g31543 not n6453 ; n6453_not
g31544 not n6525 ; n6525_not
g31545 not n8334 ; n8334_not
g31546 not n6435 ; n6435_not
g31547 not n2817 ; n2817_not
g31548 not n2835 ; n2835_not
g31549 not n2871 ; n2871_not
g31550 not n7362 ; n7362_not
g31551 not n4626 ; n4626_not
g31552 not n9316 ; n9316_not
g31553 not n7525 ; n7525_not
g31554 not n7075 ; n7075_not
g31555 not n7570 ; n7570_not
g31556 not n5770 ; n5770_not
g31557 not n7903 ; n7903_not
g31558 not n9604 ; n9604_not
g31559 not n9613 ; n9613_not
g31560 not n2485 ; n2485_not
g31561 not n7066 ; n7066_not
g31562 not n9631 ; n9631_not
g31563 not n6814 ; n6814_not
g31564 not n9361 ; n9361_not
g31565 not n7048 ; n7048_not
g31566 not n6436 ; n6436_not
g31567 not n5914 ; n5914_not
g31568 not n9910 ; n9910_not
g31569 not n6742 ; n6742_not
g31570 not n6373 ; n6373_not
g31571 not n6535 ; n6535_not
g31572 not n6355 ; n6355_not
g31573 not n8092 ; n8092_not
g31574 not n7129 ; n7129_not
g31575 not n7291 ; n7291_not
g31576 not n9622 ; n9622_not
g31577 not n7813 ; n7813_not
g31578 not n5752 ; n5752_not
g31579 not n9343 ; n9343_not
g31580 not n5716 ; n5716_not
g31581 not n7462 ; n7462_not
g31582 not n6526 ; n6526_not
g31583 not n7921 ; n7921_not
g31584 not n6517 ; n6517_not
g31585 not n6427 ; n6427_not
g31586 not n6634 ; n6634_not
g31587 not n7543 ; n7543_not
g31588 not n7507 ; n7507_not
g31589 not n7822 ; n7822_not
g31590 not n7552 ; n7552_not
g31591 not n7840 ; n7840_not
g31592 not n9352 ; n9352_not
g31593 not n6364 ; n6364_not
g31594 not n5932 ; n5932_not
g31595 not n5923 ; n5923_not
g31596 not n6706 ; n6706_not
g31597 not n5572 ; n5572_not
g31598 not n7516 ; n7516_not
g31599 not n9541 ; n9541_not
g31600 not n7057 ; n7057_not
g31601 not n7471 ; n7471_not
g31602 not n8056 ; n8056_not
g31603 not n5824 ; n5824_not
g31604 not n6472 ; n6472_not
g31605 not n6724 ; n6724_not
g31606 not n5851 ; n5851_not
g31607 not n5815 ; n5815_not
g31608 not n5743 ; n5743_not
g31609 not n9460 ; n9460_not
g31610 not n8038 ; n8038_not
g31611 not n9532 ; n9532_not
g31612 not n5842 ; n5842_not
g31613 not n6715 ; n6715_not
g31614 not n9712 ; n9712_not
g31615 not n9217 ; n9217_not
g31616 not n9730 ; n9730_not
g31617 not n6463 ; n6463_not
g31618 not n7480 ; n7480_not
g31619 not n5833 ; n5833_not
g31620 not n7930 ; n7930_not
g31621 not n9523 ; n9523_not
g31622 not n9514 ; n9514_not
g31623 not n7912 ; n7912_not
g31624 not n9424 ; n9424_not
g31625 not n8083 ; n8083_not
g31626 not n9415 ; n9415_not
g31627 not n5806 ; n5806_not
g31628 not n6382 ; n6382_not
g31629 not n6490 ; n6490_not
g31630 not n6229 ; n6229_not
g31631 not n6283 ; n6283_not
g31632 not n9406 ; n9406_not
g31633 not n9901 ; n9901_not
g31634 not n6454 ; n6454_not
g31635 not n5536 ; n5536_not
g31636 not n6418 ; n6418_not
g31637 not n6733 ; n6733_not
g31638 not n9811 ; n9811_not
g31639 not n9442 ; n9442_not
g31640 not n9802 ; n9802_not
g31641 not n8065 ; n8065_not
g31642 not n5860 ; n5860_not
g31643 not n5950 ; n5950_not
g31644 not n8074 ; n8074_not
g31645 not n7561 ; n7561_not
g31646 not n9550 ; n9550_not
g31647 not n6643 ; n6643_not
g31648 not n5941 ; n5941_not
g31649 not n6391 ; n6391_not
g31650 not n9703 ; n9703_not
g31651 not n7255 ; n7255_not
g31652 not n7363 ; n7363_not
g31653 not n7246 ; n7246_not
g31654 not n8650 ; n8650_not
g31655 not n8830 ; n8830_not
g31656 not n8821 ; n8821_not
g31657 not n8371 ; n8371_not
g31658 not n6850 ; n6850_not
g31659 not n8353 ; n8353_not
g31660 not n8812 ; n8812_not
g31661 not n7264 ; n7264_not
g31662 not n8803 ; n8803_not
g31663 not n6832 ; n6832_not
g31664 not n6166 ; n6166_not
g31665 not n7345 ; n7345_not
g31666 not n7534 ; n7534_not
g31667 not n7336 ; n7336_not
g31668 not n6175 ; n6175_not
g31669 not n8740 ; n8740_not
g31670 not n8731 ; n8731_not
g31671 not n8416 ; n8416_not
g31672 not n8407 ; n8407_not
g31673 not n8281 ; n8281_not
g31674 not n9019 ; n9019_not
g31675 not n6256 ; n6256_not
g31676 not n6157 ; n6157_not
g31677 not n7219 ; n7219_not
g31678 not n8290 ; n8290_not
g31679 not n6823 ; n6823_not
g31680 not n7381 ; n7381_not
g31681 not n8317 ; n8317_not
g31682 not n7228 ; n7228_not
g31683 not n7705 ; n7705_not
g31684 not n8335 ; n8335_not
g31685 not n7237 ; n7237_not
g31686 not n8623 ; n8623_not
g31687 not n6571 ; n6571_not
g31688 not n6247 ; n6247_not
g31689 not n8920 ; n8920_not
g31690 not n6184 ; n6184_not
g31691 not n6562 ; n6562_not
g31692 not n8344 ; n8344_not
g31693 not n8911 ; n8911_not
g31694 not n7372 ; n7372_not
g31695 not n8902 ; n8902_not
g31696 not n6922 ; n6922_not
g31697 not n8461 ; n8461_not
g31698 not n8191 ; n8191_not
g31699 not n7318 ; n7318_not
g31700 not n6913 ; n6913_not
g31701 not n8614 ; n8614_not
g31702 not n8605 ; n8605_not
g31703 not n8272 ; n8272_not
g31704 not n8551 ; n8551_not
g31705 not n8236 ; n8236_not
g31706 not n8542 ; n8542_not
g31707 not n8506 ; n8506_not
g31708 not n6904 ; n6904_not
g31709 not n8533 ; n8533_not
g31710 not n6841 ; n6841_not
g31711 not n8218 ; n8218_not
g31712 not n7723 ; n7723_not
g31713 not n7309 ; n7309_not
g31714 not n8524 ; n8524_not
g31715 not n6661 ; n6661_not
g31716 not n8515 ; n8515_not
g31717 not n7327 ; n7327_not
g31718 not n8326 ; n8326_not
g31719 not n7273 ; n7273_not
g31720 not n8722 ; n8722_not
g31721 not n8425 ; n8425_not
g31722 not n6193 ; n6193_not
g31723 not n6544 ; n6544_not
g31724 not n8713 ; n8713_not
g31725 not n8434 ; n8434_not
g31726 not n6940 ; n6940_not
g31727 not n8443 ; n8443_not
g31728 not n7282 ; n7282_not
g31729 not n8641 ; n8641_not
g31730 not n8632 ; n8632_not
g31731 not n6238 ; n6238_not
g31732 not n8452 ; n8452_not
g31733 not n6931 ; n6931_not
g31734 not n6094 ; n6094_not
g31735 not n7147 ; n7147_not
g31736 not n9226 ; n9226_not
g31737 not n6805 ; n6805_not
g31738 not n6292 ; n6292_not
g31739 not n6652 ; n6652_not
g31740 not n8137 ; n8137_not
g31741 not n7435 ; n7435_not
g31742 not n9208 ; n9208_not
g31743 not n7165 ; n7165_not
g31744 not n9190 ; n9190_not
g31745 not n7750 ; n7750_not
g31746 not n9172 ; n9172_not
g31747 not n7426 ; n7426_not
g31748 not n6607 ; n6607_not
g31749 not n8146 ; n8146_not
g31750 not n9163 ; n9163_not
g31751 not n7156 ; n7156_not
g31752 not n8155 ; n8155_not
g31753 not n7624 ; n7624_not
g31754 not n9154 ; n9154_not
g31755 not n6346 ; n6346_not
g31756 not n9325 ; n9325_not
g31757 not n7606 ; n7606_not
g31758 not n6067 ; n6067_not
g31759 not n6751 ; n6751_not
g31760 not n6337 ; n6337_not
g31761 not n9307 ; n9307_not
g31762 not n8119 ; n8119_not
g31763 not n6760 ; n6760_not
g31764 not n9253 ; n9253_not
g31765 not n9280 ; n9280_not
g31766 not n9262 ; n9262_not
g31767 not n9271 ; n9271_not
g31768 not n7453 ; n7453_not
g31769 not n6616 ; n6616_not
g31770 not n8128 ; n8128_not
g31771 not n6085 ; n6085_not
g31772 not n9244 ; n9244_not
g31773 not n7615 ; n7615_not
g31774 not n9235 ; n9235_not
g31775 not n7444 ; n7444_not
g31776 not n9082 ; n9082_not
g31777 not n9073 ; n9073_not
g31778 not n7660 ; n7660_not
g31779 not n9064 ; n9064_not
g31780 not n7408 ; n7408_not
g31781 not n9055 ; n9055_not
g31782 not n7138 ; n7138_not
g31783 not n7192 ; n7192_not
g31784 not n9046 ; n9046_not
g31785 not n8254 ; n8254_not
g31786 not n8263 ; n8263_not
g31787 not n7732 ; n7732_not
g31788 not n6265 ; n6265_not
g31789 not n7390 ; n7390_not
g31790 not n6148 ; n6148_not
g31791 not n6580 ; n6580_not
g31792 not n9028 ; n9028_not
g31793 not n8164 ; n8164_not
g31794 not n9145 ; n9145_not
g31795 not n7741 ; n7741_not
g31796 not n8173 ; n8173_not
g31797 not n8182 ; n8182_not
g31798 not n7633 ; n7633_not
g31799 not n9136 ; n9136_not
g31800 not n9127 ; n9127_not
g31801 not n7174 ; n7174_not
g31802 not n8209 ; n8209_not
g31803 not n9118 ; n9118_not
g31804 not n8029 ; n8029_not
g31805 not n7642 ; n7642_not
g31806 not n9109 ; n9109_not
g31807 not n9091 ; n9091_not
g31808 not n8227 ; n8227_not
g31809 not n4780 ; n4780_not
g31810 not n1927 ; n1927_not
g31811 not n1936 ; n1936_not
g31812 not n1873 ; n1873_not
g31813 not n4771 ; n4771_not
g31814 not n4762 ; n4762_not
g31815 not n1945 ; n1945_not
g31816 not n4753 ; n4753_not
g31817 not n4744 ; n4744_not
g31818 not n1954 ; n1954_not
g31819 not n1963 ; n1963_not
g31820 not n1981 ; n1981_not
g31821 not n1990 ; n1990_not
g31822 not n1918 ; n1918_not
g31823 not n4717 ; n4717_not
g31824 not n4690 ; n4690_not
g31825 not n1819 ; n1819_not
g31826 not n4861 ; n4861_not
g31827 not n1828 ; n1828_not
g31828 not n1837 ; n1837_not
g31829 not n4852 ; n4852_not
g31830 not n1855 ; n1855_not
g31831 not n4843 ; n4843_not
g31832 not n1864 ; n1864_not
g31833 not n4834 ; n4834_not
g31834 not n4825 ; n4825_not
g31835 not n4735 ; n4735_not
g31836 not n4816 ; n4816_not
g31837 not n1882 ; n1882_not
g31838 not n1891 ; n1891_not
g31839 not n1909 ; n1909_not
g31840 not n4663 ; n4663_not
g31841 not n4654 ; n4654_not
g31842 not n4645 ; n4645_not
g31843 not n4636 ; n4636_not
g31844 not n4627 ; n4627_not
g31845 not n2449 ; n2449_not
g31846 not n4618 ; n4618_not
g31847 not n2296 ; n2296_not
g31848 not n4357 ; n4357_not
g31849 not n4609 ; n4609_not
g31850 not n2467 ; n2467_not
g31851 not n2476 ; n2476_not
g31852 not n4591 ; n4591_not
g31853 not n2494 ; n2494_not
g31854 not n2548 ; n2548_not
g31855 not n2557 ; n2557_not
g31856 not n2566 ; n2566_not
g31857 not n2575 ; n2575_not
g31858 not n2089 ; n2089_not
g31859 not n2098 ; n2098_not
g31860 not n4681 ; n4681_not
g31861 not n2179 ; n2179_not
g31862 not n2188 ; n2188_not
g31863 not n4672 ; n4672_not
g31864 not n2278 ; n2278_not
g31865 not n2269 ; n2269_not
g31866 not n2287 ; n2287_not
g31867 not n2359 ; n2359_not
g31868 not n2368 ; n2368_not
g31869 not n2377 ; n2377_not
g31870 not n2386 ; n2386_not
g31871 not n5437 ; n5437_not
g31872 not n5428 ; n5428_not
g31873 not n5419 ; n5419_not
g31874 not n5392 ; n5392_not
g31875 not n5248 ; n5248_not
g31876 not n5383 ; n5383_not
g31877 not n5374 ; n5374_not
g31878 not n5365 ; n5365_not
g31879 not n5356 ; n5356_not
g31880 not n5347 ; n5347_not
g31881 not n5329 ; n5329_not
g31882 not n5293 ; n5293_not
g31883 not n5284 ; n5284_not
g31884 not n5275 ; n5275_not
g31885 not n1594 ; n1594_not
g31886 not n5581 ; n5581_not
g31887 not n5590 ; n5590_not
g31888 not n1486 ; n1486_not
g31889 not n1549 ; n1549_not
g31890 not n5563 ; n5563_not
g31891 not n1567 ; n1567_not
g31892 not n5554 ; n5554_not
g31893 not n5545 ; n5545_not
g31894 not n5527 ; n5527_not
g31895 not n5509 ; n5509_not
g31896 not n1459 ; n1459_not
g31897 not n1576 ; n1576_not
g31898 not n5491 ; n5491_not
g31899 not n5482 ; n5482_not
g31900 not n5473 ; n5473_not
g31901 not n5455 ; n5455_not
g31902 not n5446 ; n5446_not
g31903 not n1684 ; n1684_not
g31904 not n1693 ; n1693_not
g31905 not n4960 ; n4960_not
g31906 not n4951 ; n4951_not
g31907 not n1729 ; n1729_not
g31908 not n1747 ; n1747_not
g31909 not n4933 ; n4933_not
g31910 not n1756 ; n1756_not
g31911 not n1765 ; n1765_not
g31912 not n1774 ; n1774_not
g31913 not n4924 ; n4924_not
g31914 not n1783 ; n1783_not
g31915 not n4906 ; n4906_not
g31916 not n1792 ; n1792_not
g31917 not n4870 ; n4870_not
g31918 not n5257 ; n5257_not
g31919 not n5239 ; n5239_not
g31920 not n1639 ; n1639_not
g31921 not n1648 ; n1648_not
g31922 not n5194 ; n5194_not
g31923 not n1657 ; n1657_not
g31924 not n5185 ; n5185_not
g31925 not n5176 ; n5176_not
g31926 not n5167 ; n5167_not
g31927 not n5158 ; n5158_not
g31928 not n5149 ; n5149_not
g31929 not n5095 ; n5095_not
g31930 not n5086 ; n5086_not
g31931 not n5077 ; n5077_not
g31932 not n5068 ; n5068_not
g31933 not n1666 ; n1666_not
g31934 not n5059 ; n5059_not
g31935 not n2917 ; n2917_not
g31936 not n3754 ; n3754_not
g31937 not n3745 ; n3745_not
g31938 not n2926 ; n2926_not
g31939 not n3736 ; n3736_not
g31940 not n3727 ; n3727_not
g31941 not n2656 ; n2656_not
g31942 not n2935 ; n2935_not
g31943 not n3718 ; n3718_not
g31944 not n2944 ; n2944_not
g31945 not n2953 ; n2953_not
g31946 not n2962 ; n2962_not
g31947 not n2782 ; n2782_not
g31948 not n3709 ; n3709_not
g31949 not n2971 ; n2971_not
g31950 not n3691 ; n3691_not
g31951 not n2980 ; n2980_not
g31952 not n2809 ; n2809_not
g31953 not n3637 ; n3637_not
g31954 not n3628 ; n3628_not
g31955 not n3835 ; n3835_not
g31956 not n3826 ; n3826_not
g31957 not n3808 ; n3808_not
g31958 not n2863 ; n2863_not
g31959 not n3790 ; n3790_not
g31960 not n2881 ; n2881_not
g31961 not n2890 ; n2890_not
g31962 not n2872 ; n2872_not
g31963 not n3781 ; n3781_not
g31964 not n2908 ; n2908_not
g31965 not n3772 ; n3772_not
g31966 not n3763 ; n3763_not
g31967 not n3367 ; n3367_not
g31968 not n3187 ; n3187_not
g31969 not n3619 ; n3619_not
g31970 not n3385 ; n3385_not
g31971 not n3394 ; n3394_not
g31972 not n3592 ; n3592_not
g31973 not n3439 ; n3439_not
g31974 not n3448 ; n3448_not
g31975 not n3457 ; n3457_not
g31976 not n3583 ; n3583_not
g31977 not n3475 ; n3475_not
g31978 not n3493 ; n3493_not
g31979 not n3538 ; n3538_not
g31980 not n3529 ; n3529_not
g31981 not n3547 ; n3547_not
g31982 not n3556 ; n3556_not
g31983 not n3574 ; n3574_not
g31984 not n3682 ; n3682_not
g31985 not n3673 ; n3673_not
g31986 not n3088 ; n3088_not
g31987 not n3178 ; n3178_not
g31988 not n3196 ; n3196_not
g31989 not n3259 ; n3259_not
g31990 not n3268 ; n3268_not
g31991 not n3664 ; n3664_not
g31992 not n3655 ; n3655_not
g31993 not n3277 ; n3277_not
g31994 not n3286 ; n3286_not
g31995 not n3295 ; n3295_not
g31996 not n3646 ; n3646_not
g31997 not n3358 ; n3358_not
g31998 not n4447 ; n4447_not
g31999 not n4438 ; n4438_not
g32000 not n4186 ; n4186_not
g32001 not n4429 ; n4429_not
g32002 not n4393 ; n4393_not
g32003 not n4384 ; n4384_not
g32004 not n4375 ; n4375_not
g32005 not n4366 ; n4366_not
g32006 not n4348 ; n4348_not
g32007 not n4339 ; n4339_not
g32008 not n4294 ; n4294_not
g32009 not n4285 ; n4285_not
g32010 not n4276 ; n4276_not
g32011 not n4267 ; n4267_not
g32012 not n4249 ; n4249_not
g32013 not n4195 ; n4195_not
g32014 not n2584 ; n2584_not
g32015 not n2593 ; n2593_not
g32016 not n2629 ; n2629_not
g32017 not n2638 ; n2638_not
g32018 not n2647 ; n2647_not
g32019 not n4528 ; n4528_not
g32020 not n4564 ; n4564_not
g32021 not n4573 ; n4573_not
g32022 not n4555 ; n4555_not
g32023 not n4546 ; n4546_not
g32024 not n4537 ; n4537_not
g32025 not n4519 ; n4519_not
g32026 not n4492 ; n4492_not
g32027 not n2665 ; n2665_not
g32028 not n4483 ; n4483_not
g32029 not n2674 ; n2674_not
g32030 not n4474 ; n4474_not
g32031 not n4465 ; n4465_not
g32032 not n4456 ; n4456_not
g32033 not n2773 ; n2773_not
g32034 not n3934 ; n3934_not
g32035 not n3925 ; n3925_not
g32036 not n3916 ; n3916_not
g32037 not n3907 ; n3907_not
g32038 not n2791 ; n2791_not
g32039 not n3871 ; n3871_not
g32040 not n2818 ; n2818_not
g32041 not n2827 ; n2827_not
g32042 not n2836 ; n2836_not
g32043 not n3862 ; n3862_not
g32044 not n2845 ; n2845_not
g32045 not n3853 ; n3853_not
g32046 not n3844 ; n3844_not
g32047 not n2683 ; n2683_not
g32048 not n4168 ; n4168_not
g32049 not n4177 ; n4177_not
g32050 not n2692 ; n2692_not
g32051 not n4159 ; n4159_not
g32052 not n4087 ; n4087_not
g32053 not n4078 ; n4078_not
g32054 not n4069 ; n4069_not
g32055 not n3970 ; n3970_not
g32056 not n2719 ; n2719_not
g32057 not n2728 ; n2728_not
g32058 not n2737 ; n2737_not
g32059 not n2746 ; n2746_not
g32060 not n2755 ; n2755_not
g32061 not n1288 ; n1288_not
g32062 not n5707 ; n5707_not
g32063 not n5680 ; n5680_not
g32064 not n1396 ; n1396_not
g32065 not n1198 ; n1198_not
g32066 not n5635 ; n5635_not
g32067 not n1468 ; n1468_not
g32068 not n1378 ; n1378_not
g32069 not n5662 ; n5662_not
g32070 not n1189 ; n1189_not
g32071 not n1369 ; n1369_not
g32072 not n1279 ; n1279_not
g32073 not n5644 ; n5644_not
g32074 not n5608 ; n5608_not
g32075 not n5653 ; n5653_not
g32076 not n1387 ; n1387_not
g32077 not n1477 ; n1477_not
g32078 not n5671 ; n5671_not
g32079 not n1495 ; n1495_not
g32080 not n5617 ; n5617_not
g32081 not n5725 ; n5725_not
g32082 not n5626 ; n5626_not
g32083 not n1099 ; n1099_not
g32084 not n2099 ; n2099_not
g32085 not n6716 ; n6716_not
g32086 not n9074 ; n9074_not
g32087 not n6734 ; n6734_not
g32088 not n8219 ; n8219_not
g32089 not n6419 ; n6419_not
g32090 not n3485 ; n3485_not
g32091 not n2837 ; n2837_not
g32092 not n5654 ; n5654_not
g32093 not n9065 ; n9065_not
g32094 not n2972 ; n2972_not
g32095 not n6725 ; n6725_not
g32096 not n7634 ; n7634_not
g32097 not n1973 ; n1973_not
g32098 not n9119 ; n9119_not
g32099 not n3476 ; n3476_not
g32100 not n1982 ; n1982_not
g32101 not n8192 ; n8192_not
g32102 not n9056 ; n9056_not
g32103 not n1991 ; n1991_not
g32104 not n6680 ; n6680_not
g32105 not n4664 ; n4664_not
g32106 not n7625 ; n7625_not
g32107 not n3683 ; n3683_not
g32108 not n2981 ; n2981_not
g32109 not n9092 ; n9092_not
g32110 not n1793 ; n1793_not
g32111 not n7616 ; n7616_not
g32112 not n5906 ; n5906_not
g32113 not n5771 ; n5771_not
g32114 not n4718 ; n4718_not
g32115 not n4709 ; n4709_not
g32116 not n6707 ; n6707_not
g32117 not n9083 ; n9083_not
g32118 not n3692 ; n3692_not
g32119 not n7607 ; n7607_not
g32120 not n4691 ; n4691_not
g32121 not n8633 ; n8633_not
g32122 not n9713 ; n9713_not
g32123 not n8606 ; n8606_not
g32124 not n8930 ; n8930_not
g32125 not n7571 ; n7571_not
g32126 not n8921 ; n8921_not
g32127 not n6806 ; n6806_not
g32128 not n4655 ; n4655_not
g32129 not n3719 ; n3719_not
g32130 not n4646 ; n4646_not
g32131 not n2927 ; n2927_not
g32132 not n6815 ; n6815_not
g32133 not n4637 ; n4637_not
g32134 not n9722 ; n9722_not
g32135 not n4628 ; n4628_not
g32136 not n5663 ; n5663_not
g32137 not n6824 ; n6824_not
g32138 not n8912 ; n8912_not
g32139 not n8255 ; n8255_not
g32140 not n6833 ; n6833_not
g32141 not n7562 ; n7562_not
g32142 not n2459 ; n2459_not
g32143 not n9047 ; n9047_not
g32144 not n6743 ; n6743_not
g32145 not n2189 ; n2189_not
g32146 not n4673 ; n4673_not
g32147 not n2963 ; n2963_not
g32148 not n1397 ; n1397_not
g32149 not n6446 ; n6446_not
g32150 not n6752 ; n6752_not
g32151 not n2279 ; n2279_not
g32152 not n2954 ; n2954_not
g32153 not n9029 ; n9029_not
g32154 not n2297 ; n2297_not
g32155 not n6770 ; n6770_not
g32156 not n1298 ; n1298_not
g32157 not n2378 ; n2378_not
g32158 not n8237 ; n8237_not
g32159 not n2369 ; n2369_not
g32160 not n2387 ; n2387_not
g32161 not n2396 ; n2396_not
g32162 not n7580 ; n7580_not
g32163 not n2945 ; n2945_not
g32164 not n8066 ; n8066_not
g32165 not n1856 ; n1856_not
g32166 not n3197 ; n3197_not
g32167 not n4844 ; n4844_not
g32168 not n9227 ; n9227_not
g32169 not n3188 ; n3188_not
g32170 not n4835 ; n4835_not
g32171 not n9650 ; n9650_not
g32172 not n8129 ; n8129_not
g32173 not n9902 ; n9902_not
g32174 not n6509 ; n6509_not
g32175 not n5717 ; n5717_not
g32176 not n4826 ; n4826_not
g32177 not n3179 ; n3179_not
g32178 not n6518 ; n6518_not
g32179 not n9641 ; n9641_not
g32180 not n4817 ; n4817_not
g32181 not n4583 ; n4583_not
g32182 not n5924 ; n5924_not
g32183 not n3089 ; n3089_not
g32184 not n1874 ; n1874_not
g32185 not n5483 ; n5483_not
g32186 not n1883 ; n1883_not
g32187 not n9209 ; n9209_not
g32188 not n6536 ; n6536_not
g32189 not n5708 ; n5708_not
g32190 not n6257 ; n6257_not
g32191 not n4871 ; n4871_not
g32192 not n1757 ; n1757_not
g32193 not n6455 ; n6455_not
g32194 not n9263 ; n9263_not
g32195 not n9821 ; n9821_not
g32196 not n3656 ; n3656_not
g32197 not n4862 ; n4862_not
g32198 not n5933 ; n5933_not
g32199 not n3269 ; n3269_not
g32200 not n6464 ; n6464_not
g32201 not n9254 ; n9254_not
g32202 not n1829 ; n1829_not
g32203 not n7706 ; n7706_not
g32204 not n4853 ; n4853_not
g32205 not n6473 ; n6473_not
g32206 not n5762 ; n5762_not
g32207 not n9245 ; n9245_not
g32208 not n3665 ; n3665_not
g32209 not n1847 ; n1847_not
g32210 not n9236 ; n9236_not
g32211 not n6491 ; n6491_not
g32212 not n8183 ; n8183_not
g32213 not n6572 ; n6572_not
g32214 not n8804 ; n8804_not
g32215 not n4763 ; n4763_not
g32216 not n6329 ; n6329_not
g32217 not n6617 ; n6617_not
g32218 not n9146 ; n9146_not
g32219 not n7652 ; n7652_not
g32220 not n1946 ; n1946_not
g32221 not n4754 ; n4754_not
g32222 not n7643 ; n7643_not
g32223 not n4745 ; n4745_not
g32224 not n3674 ; n3674_not
g32225 not n1955 ; n1955_not
g32226 not n4736 ; n4736_not
g32227 not n9137 ; n9137_not
g32228 not n1964 ; n1964_not
g32229 not n6653 ; n6653_not
g32230 not n9128 ; n9128_not
g32231 not n4727 ; n4727_not
g32232 not n6662 ; n6662_not
g32233 not n1892 ; n1892_not
g32234 not n6545 ; n6545_not
g32235 not n6554 ; n6554_not
g32236 not n8147 ; n8147_not
g32237 not n2891 ; n2891_not
g32238 not n6563 ; n6563_not
g32239 not n9191 ; n9191_not
g32240 not n8156 ; n8156_not
g32241 not n8165 ; n8165_not
g32242 not n9173 ; n9173_not
g32243 not n1775 ; n1775_not
g32244 not n6581 ; n6581_not
g32245 not n5636 ; n5636_not
g32246 not n4781 ; n4781_not
g32247 not n8822 ; n8822_not
g32248 not n9164 ; n9164_not
g32249 not n7661 ; n7661_not
g32250 not n1919 ; n1919_not
g32251 not n1937 ; n1937_not
g32252 not n9155 ; n9155_not
g32253 not n8174 ; n8174_not
g32254 not n4772 ; n4772_not
g32255 not n6608 ; n6608_not
g32256 not n5915 ; n5915_not
g32257 not n4259 ; n4259_not
g32258 not n1289 ; n1289_not
g32259 not n8543 ; n8543_not
g32260 not n7148 ; n7148_not
g32261 not n2558 ; n2558_not
g32262 not n8534 ; n8534_not
g32263 not n3854 ; n3854_not
g32264 not n6914 ; n6914_not
g32265 not n4196 ; n4196_not
g32266 not n8381 ; n8381_not
g32267 not n7157 ; n7157_not
g32268 not n4187 ; n4187_not
g32269 not n7166 ; n7166_not
g32270 not n5834 ; n5834_not
g32271 not n4178 ; n4178_not
g32272 not n4169 ; n4169_not
g32273 not n8390 ; n8390_not
g32274 not n7175 ; n7175_not
g32275 not n7391 ; n7391_not
g32276 not n3863 ; n3863_not
g32277 not n7184 ; n7184_not
g32278 not n2693 ; n2693_not
g32279 not n4088 ; n4088_not
g32280 not n7193 ; n7193_not
g32281 not n4079 ; n4079_not
g32282 not n7382 ; n7382_not
g32283 not n8525 ; n8525_not
g32284 not n3827 ; n3827_not
g32285 not n7085 ; n7085_not
g32286 not n4385 ; n4385_not
g32287 not n5843 ; n5843_not
g32288 not n7094 ; n7094_not
g32289 not n7427 ; n7427_not
g32290 not n4376 ; n4376_not
g32291 not n8372 ; n8372_not
g32292 not n4367 ; n4367_not
g32293 not n9533 ; n9533_not
g32294 not n4349 ; n4349_not
g32295 not n5672 ; n5672_not
g32296 not n4277 ; n4277_not
g32297 not n8561 ; n8561_not
g32298 not n7418 ; n7418_not
g32299 not n4295 ; n4295_not
g32300 not n8552 ; n8552_not
g32301 not n2675 ; n2675_not
g32302 not n4286 ; n4286_not
g32303 not n3845 ; n3845_not
g32304 not n2846 ; n2846_not
g32305 not n7409 ; n7409_not
g32306 not n9812 ; n9812_not
g32307 not n4268 ; n4268_not
g32308 not n7139 ; n7139_not
g32309 not n3953 ; n3953_not
g32310 not n8462 ; n8462_not
g32311 not n3872 ; n3872_not
g32312 not n8453 ; n8453_not
g32313 not n8327 ; n8327_not
g32314 not n7283 ; n7283_not
g32315 not n7346 ; n7346_not
g32316 not n2765 ; n2765_not
g32317 not n8444 ; n8444_not
g32318 not n3881 ; n3881_not
g32319 not n3944 ; n3944_not
g32320 not n2774 ; n2774_not
g32321 not n7292 ; n7292_not
g32322 not n3935 ; n3935_not
g32323 not n3836 ; n3836_not
g32324 not n2792 ; n2792_not
g32325 not n3926 ; n3926_not
g32326 not n9830 ; n9830_not
g32327 not n5816 ; n5816_not
g32328 not n7337 ; n7337_not
g32329 not n7319 ; n7319_not
g32330 not n8435 ; n8435_not
g32331 not n8426 ; n8426_not
g32332 not n3890 ; n3890_not
g32333 not n7328 ; n7328_not
g32334 not n2549 ; n2549_not
g32335 not n5681 ; n5681_not
g32336 not n5825 ; n5825_not
g32337 not n2729 ; n2729_not
g32338 not n2738 ; n2738_not
g32339 not n2828 ; n2828_not
g32340 not n8507 ; n8507_not
g32341 not n7229 ; n7229_not
g32342 not n2819 ; n2819_not
g32343 not n3980 ; n3980_not
g32344 not n3764 ; n3764_not
g32345 not n2756 ; n2756_not
g32346 not n2747 ; n2747_not
g32347 not n3971 ; n3971_not
g32348 not n7364 ; n7364_not
g32349 not n7247 ; n7247_not
g32350 not n8408 ; n8408_not
g32351 not n8480 ; n8480_not
g32352 not n7256 ; n7256_not
g32353 not n8471 ; n8471_not
g32354 not n8417 ; n8417_not
g32355 not n7355 ; n7355_not
g32356 not n7265 ; n7265_not
g32357 not n6932 ; n6932_not
g32358 not n8741 ; n8741_not
g32359 not n2909 ; n2909_not
g32360 not n3773 ; n3773_not
g32361 not n8723 ; n8723_not
g32362 not n6950 ; n6950_not
g32363 not n6941 ; n6941_not
g32364 not n9911 ; n9911_not
g32365 not n8291 ; n8291_not
g32366 not n9740 ; n9740_not
g32367 not n2576 ; n2576_not
g32368 not n2585 ; n2585_not
g32369 not n7490 ; n7490_not
g32370 not n8318 ; n8318_not
g32371 not n8660 ; n8660_not
g32372 not n8651 ; n8651_not
g32373 not n3782 ; n3782_not
g32374 not n2882 ; n2882_not
g32375 not n7472 ; n7472_not
g32376 not n7481 ; n7481_not
g32377 not n7553 ; n7553_not
g32378 not n3728 ; n3728_not
g32379 not n6860 ; n6860_not
g32380 not n8840 ; n8840_not
g32381 not n7544 ; n7544_not
g32382 not n3737 ; n3737_not
g32383 not n8831 ; n8831_not
g32384 not n2468 ; n2468_not
g32385 not n8813 ; n8813_not
g32386 not n7535 ; n7535_not
g32387 not n2486 ; n2486_not
g32388 not n4592 ; n4592_not
g32389 not n2918 ; n2918_not
g32390 not n9353 ; n9353_not
g32391 not n7526 ; n7526_not
g32392 not n3755 ; n3755_not
g32393 not n8273 ; n8273_not
g32394 not n6923 ; n6923_not
g32395 not n8750 ; n8750_not
g32396 not n2495 ; n2495_not
g32397 not n7454 ; n7454_not
g32398 not n4493 ; n4493_not
g32399 not n2657 ; n2657_not
g32400 not n8354 ; n8354_not
g32401 not n2666 ; n2666_not
g32402 not n8363 ; n8363_not
g32403 not n3584 ; n3584_not
g32404 not n7049 ; n7049_not
g32405 not n7445 ; n7445_not
g32406 not n4475 ; n4475_not
g32407 not n3809 ; n3809_not
g32408 not n9704 ; n9704_not
g32409 not n7058 ; n7058_not
g32410 not n4457 ; n4457_not
g32411 not n4448 ; n4448_not
g32412 not n2855 ; n2855_not
g32413 not n7067 ; n7067_not
g32414 not n9803 ; n9803_not
g32415 not n3818 ; n3818_not
g32416 not n7076 ; n7076_not
g32417 not n4394 ; n4394_not
g32418 not n1199 ; n1199_not
g32419 not n8570 ; n8570_not
g32420 not n5870 ; n5870_not
g32421 not n2594 ; n2594_not
g32422 not n6851 ; n6851_not
g32423 not n2873 ; n2873_not
g32424 not n8624 ; n8624_not
g32425 not n2639 ; n2639_not
g32426 not n3575 ; n3575_not
g32427 not n8336 ; n8336_not
g32428 not n2648 ; n2648_not
g32429 not n8615 ; n8615_not
g32430 not n4574 ; n4574_not
g32431 not n4565 ; n4565_not
g32432 not n4529 ; n4529_not
g32433 not n3791 ; n3791_not
g32434 not n4556 ; n4556_not
g32435 not n7463 ; n7463_not
g32436 not n5861 ; n5861_not
g32437 not n4547 ; n4547_not
g32438 not n4538 ; n4538_not
g32439 not n7436 ; n7436_not
g32440 not n2864 ; n2864_not
g32441 not n5159 ; n5159_not
g32442 not n4961 ; n4961_not
g32443 not n6239 ; n6239_not
g32444 not n9416 ; n9416_not
g32445 not n3449 ; n3449_not
g32446 not n3593 ; n3593_not
g32447 not n5096 ; n5096_not
g32448 not n6248 ; n6248_not
g32449 not n5960 ; n5960_not
g32450 not n5087 ; n5087_not
g32451 not n5078 ; n5078_not
g32452 not n6167 ; n6167_not
g32453 not n5726 ; n5726_not
g32454 not n6266 ; n6266_not
g32455 not n1658 ; n1658_not
g32456 not n5069 ; n5069_not
g32457 not n1388 ; n1388_not
g32458 not n9920 ; n9920_not
g32459 not n9434 ; n9434_not
g32460 not n5258 ; n5258_not
g32461 not n8039 ; n8039_not
g32462 not n5249 ; n5249_not
g32463 not n9614 ; n9614_not
g32464 not n5168 ; n5168_not
g32465 not n9425 ; n9425_not
g32466 not n5177 ; n5177_not
g32467 not n5951 ; n5951_not
g32468 not n5195 ; n5195_not
g32469 not n1649 ; n1649_not
g32470 not n9623 ; n9623_not
g32471 not n3467 ; n3467_not
g32472 not n5186 ; n5186_not
g32473 not n3458 ; n3458_not
g32474 not n7814 ; n7814_not
g32475 not n3395 ; n3395_not
g32476 not n1694 ; n1694_not
g32477 not n3386 ; n3386_not
g32478 not n4970 ; n4970_not
g32479 not n6338 ; n6338_not
g32480 not n8084 ; n8084_not
g32481 not n9344 ; n9344_not
g32482 not n3377 ; n3377_not
g32483 not n6347 ; n6347_not
g32484 not n4952 ; n4952_not
g32485 not n8093 ; n8093_not
g32486 not n9335 ; n9335_not
g32487 not n6356 ; n6356_not
g32488 not n6284 ; n6284_not
g32489 not n5447 ; n5447_not
g32490 not n5744 ; n5744_not
g32491 not n9407 ; n9407_not
g32492 not n1667 ; n1667_not
g32493 not n7841 ; n7841_not
g32494 not n1676 ; n1676_not
g32495 not n8057 ; n8057_not
g32496 not n3296 ; n3296_not
g32497 not n1685 ; n1685_not
g32498 not n6293 ; n6293_not
g32499 not n6095 ; n6095_not
g32500 not n9632 ; n9632_not
g32501 not n5555 ; n5555_not
g32502 not n7823 ; n7823_not
g32503 not n9380 ; n9380_not
g32504 not n8075 ; n8075_not
g32505 not n9371 ; n9371_not
g32506 not n9362 ; n9362_not
g32507 not n5546 ; n5546_not
g32508 not n9560 ; n9560_not
g32509 not n7931 ; n7931_not
g32510 not n6068 ; n6068_not
g32511 not n1568 ; n1568_not
g32512 not n5609 ; n5609_not
g32513 not n7940 ; n7940_not
g32514 not n1577 ; n1577_not
g32515 not n3368 ; n3368_not
g32516 not n5492 ; n5492_not
g32517 not n6086 ; n6086_not
g32518 not n5348 ; n5348_not
g32519 not n5357 ; n5357_not
g32520 not n1586 ; n1586_not
g32521 not n5474 ; n5474_not
g32522 not n3557 ; n3557_not
g32523 not n5465 ; n5465_not
g32524 not n9551 ; n9551_not
g32525 not n5591 ; n5591_not
g32526 not n9542 ; n9542_not
g32527 not n7904 ; n7904_not
g32528 not n5582 ; n5582_not
g32529 not n7913 ; n7913_not
g32530 not n5573 ; n5573_not
g32531 not n7733 ; n7733_not
g32532 not n9524 ; n9524_not
g32533 not n5564 ; n5564_not
g32534 not n7922 ; n7922_not
g32535 not n3566 ; n3566_not
g32536 not n9515 ; n9515_not
g32537 not n5339 ; n5339_not
g32538 not n5285 ; n5285_not
g32539 not n9443 ; n9443_not
g32540 not n1469 ; n1469_not
g32541 not n6176 ; n6176_not
g32542 not n1595 ; n1595_not
g32543 not n7832 ; n7832_not
g32544 not n6185 ; n6185_not
g32545 not n5267 ; n5267_not
g32546 not n5429 ; n5429_not
g32547 not n5456 ; n5456_not
g32548 not n5438 ; n5438_not
g32549 not n9290 ; n9290_not
g32550 not n1496 ; n1496_not
g32551 not n3548 ; n3548_not
g32552 not n3539 ; n3539_not
g32553 not n5393 ; n5393_not
g32554 not n1487 ; n1487_not
g32555 not n9605 ; n9605_not
g32556 not n5780 ; n5780_not
g32557 not n5384 ; n5384_not
g32558 not n9461 ; n9461_not
g32559 not n5375 ; n5375_not
g32560 not n3494 ; n3494_not
g32561 not n7760 ; n7760_not
g32562 not n5366 ; n5366_not
g32563 not n9308 ; n9308_not
g32564 not n9281 ; n9281_not
g32565 not n4907 ; n4907_not
g32566 not n4682 ; n4682_not
g32567 not n9317 ; n9317_not
g32568 not n3287 ; n3287_not
g32569 not n9326 ; n9326_not
g32570 not n3359 ; n3359_not
g32571 not n6428 ; n6428_not
g32572 not n7742 ; n7742_not
g32573 not n6437 ; n6437_not
g32574 not n7751 ; n7751_not
g32575 not n9272 ; n9272_not
g32576 not n5753 ; n5753_not
g32577 not n4925 ; n4925_not
g32578 not n4934 ; n4934_not
g32579 not n3629 ; n3629_not
g32580 not n3647 ; n3647_not
g32581 not n3278 ; n3278_not
g32582 not n5618 ; n5618_not
g32583 not n6374 ; n6374_not
g32584 not n6392 ; n6392_not
g32585 not n7724 ; n7724_not
g32586 not n5942 ; n5942_not
g32587 not n1748 ; n1748_not
g32588 not n4916 ; n4916_not
g32589 not n1784 ; n1784_not
g32590 not n5627 ; n5627_not
g32591 not n7059 ; n7059_not
g32592 not n4278 ; n4278_not
g32593 not n5529 ; n5529_not
g32594 not n9606 ; n9606_not
g32595 not n9129 ; n9129_not
g32596 not n2856 ; n2856_not
g32597 not n7419 ; n7419_not
g32598 not n7095 ; n7095_not
g32599 not n7860 ; n7860_not
g32600 not n3549 ; n3549_not
g32601 not n9804 ; n9804_not
g32602 not n5448 ; n5448_not
g32603 not n3783 ; n3783_not
g32604 not n5385 ; n5385_not
g32605 not n5673 ; n5673_not
g32606 not n4890 ; n4890_not
g32607 not n7068 ; n7068_not
g32608 not n1776 ; n1776_not
g32609 not n8553 ; n8553_not
g32610 not n4476 ; n4476_not
g32611 not n7725 ; n7725_not
g32612 not n3198 ; n3198_not
g32613 not n9705 ; n9705_not
g32614 not n5754 ; n5754_not
g32615 not n3495 ; n3495_not
g32616 not n8562 ; n8562_not
g32617 not n4467 ; n4467_not
g32618 not n1857 ; n1857_not
g32619 not n5376 ; n5376_not
g32620 not n1587 ; n1587_not
g32621 not n3648 ; n3648_not
g32622 not n4296 ; n4296_not
g32623 not n1848 ; n1848_not
g32624 not n7851 ; n7851_not
g32625 not n4368 ; n4368_not
g32626 not n1794 ; n1794_not
g32627 not n9174 ; n9174_not
g32628 not n8571 ; n8571_not
g32629 not n2676 ; n2676_not
g32630 not n9471 ; n9471_not
g32631 not n6492 ; n6492_not
g32632 not n3828 ; n3828_not
g32633 not n4386 ; n4386_not
g32634 not n9552 ; n9552_not
g32635 not n5736 ; n5736_not
g32636 not n7428 ; n7428_not
g32637 not n5844 ; n5844_not
g32638 not n7923 ; n7923_not
g32639 not n6483 ; n6483_not
g32640 not n9291 ; n9291_not
g32641 not n9462 ; n9462_not
g32642 not n5727 ; n5727_not
g32643 not n2847 ; n2847_not
g32644 not n8580 ; n8580_not
g32645 not n9480 ; n9480_not
g32646 not n3819 ; n3819_not
g32647 not n7932 ; n7932_not
g32648 not n7077 ; n7077_not
g32649 not n4359 ; n4359_not
g32650 not n5763 ; n5763_not
g32651 not n4395 ; n4395_not
g32652 not n3738 ; n3738_not
g32653 not n8670 ; n8670_not
g32654 not n5268 ; n5268_not
g32655 not n8490 ; n8490_not
g32656 not n7833 ; n7833_not
g32657 not n8652 ; n8652_not
g32658 not n1596 ; n1596_not
g32659 not n4827 ; n4827_not
g32660 not n7482 ; n7482_not
g32661 not n9219 ; n9219_not
g32662 not n8634 ; n8634_not
g32663 not n6177 ; n6177_not
g32664 not n2595 ; n2595_not
g32665 not n4692 ; n4692_not
g32666 not n2874 ; n2874_not
g32667 not n4908 ; n4908_not
g32668 not n7473 ; n7473_not
g32669 not n4836 ; n4836_not
g32670 not n5286 ; n5286_not
g32671 not n6942 ; n6942_not
g32672 not n7509 ; n7509_not
g32673 not n9435 ; n9435_not
g32674 not n2559 ; n2559_not
g32675 not n3774 ; n3774_not
g32676 not n3189 ; n3189_not
g32677 not n6951 ; n6951_not
g32678 not n4917 ; n4917_not
g32679 not n5925 ; n5925_not
g32680 not n5790 ; n5790_not
g32681 not n7491 ; n7491_not
g32682 not n3558 ; n3558_not
g32683 not n8292 ; n8292_not
g32684 not n8706 ; n8706_not
g32685 not n6960 ; n6960_not
g32686 not n7824 ; n7824_not
g32687 not n2577 ; n2577_not
g32688 not n3468 ; n3468_not
g32689 not n9741 ; n9741_not
g32690 not n8463 ; n8463_not
g32691 not n6186 ; n6186_not
g32692 not n2892 ; n2892_not
g32693 not n4539 ; n4539_not
g32694 not n6825 ; n6825_not
g32695 not n1785 ; n1785_not
g32696 not n7842 ; n7842_not
g32697 not n5349 ; n5349_not
g32698 not n5259 ; n5259_not
g32699 not n7437 ; n7437_not
g32700 not n8607 ; n8607_not
g32701 not n5079 ; n5079_not
g32702 not n2658 ; n2658_not
g32703 not n7455 ; n7455_not
g32704 not n9228 ; n9228_not
g32705 not n4494 ; n4494_not
g32706 not n3486 ; n3486_not
g32707 not n8355 ; n8355_not
g32708 not n5367 ; n5367_not
g32709 not n9651 ; n9651_not
g32710 not n9444 ; n9444_not
g32711 not n8616 ; n8616_not
g32712 not n3477 ; n3477_not
g32713 not n6168 ; n6168_not
g32714 not n4575 ; n4575_not
g32715 not n8337 ; n8337_not
g32716 not n2649 ; n2649_not
g32717 not n1398 ; n1398_not
g32718 not n4566 ; n4566_not
g32719 not n4557 ; n4557_not
g32720 not n5934 ; n5934_not
g32721 not n4719 ; n4719_not
g32722 not n9453 ; n9453_not
g32723 not n5862 ; n5862_not
g32724 not n4548 ; n4548_not
g32725 not n3792 ; n3792_not
g32726 not n1488 ; n1488_not
g32727 not n7248 ; n7248_not
g32728 not n8481 ; n8481_not
g32729 not n9831 ; n9831_not
g32730 not n6438 ; n6438_not
g32731 not n7257 ; n7257_not
g32732 not n9561 ; n9561_not
g32733 not n8472 ; n8472_not
g32734 not n3963 ; n3963_not
g32735 not n8175 ; n8175_not
g32736 not n7356 ; n7356_not
g32737 not n3954 ; n3954_not
g32738 not n5565 ; n5565_not
g32739 not n7266 ; n7266_not
g32740 not n8418 ; n8418_not
g32741 not n5556 ; n5556_not
g32742 not n9264 ; n9264_not
g32743 not n2766 ; n2766_not
g32744 not n7086 ; n7086_not
g32745 not n3990 ; n3990_not
g32746 not n2667 ; n2667_not
g32747 not n9570 ; n9570_not
g32748 not n7707 ; n7707_not
g32749 not n5547 ; n5547_not
g32750 not n2748 ; n2748_not
g32751 not n3981 ; n3981_not
g32752 not n1569 ; n1569_not
g32753 not n9840 ; n9840_not
g32754 not n6465 ; n6465_not
g32755 not n8409 ; n8409_not
g32756 not n7239 ; n7239_not
g32757 not n7365 ; n7365_not
g32758 not n2757 ; n2757_not
g32759 not n3972 ; n3972_not
g32760 not n5457 ; n5457_not
g32761 not n9516 ; n9516_not
g32762 not n5583 ; n5583_not
g32763 not n2793 ; n2793_not
g32764 not n3927 ; n3927_not
g32765 not n3837 ; n3837_not
g32766 not n1758 ; n1758_not
g32767 not n9642 ; n9642_not
g32768 not n9822 ; n9822_not
g32769 not n7716 ; n7716_not
g32770 not n7338 ; n7338_not
g32771 not n3909 ; n3909_not
g32772 not n9543 ; n9543_not
g32773 not n7905 ; n7905_not
g32774 not n6447 ; n6447_not
g32775 not n2784 ; n2784_not
g32776 not n5592 ; n5592_not
g32777 not n8427 ; n8427_not
g32778 not n7329 ; n7329_not
g32779 not n3891 ; n3891_not
g32780 not n3657 ; n3657_not
g32781 not n8454 ; n8454_not
g32782 not n5484 ; n5484_not
g32783 not n7734 ; n7734_not
g32784 not n3945 ; n3945_not
g32785 not n7347 ; n7347_not
g32786 not n4863 ; n4863_not
g32787 not n7284 ; n7284_not
g32788 not n5835 ; n5835_not
g32789 not n8445 ; n8445_not
g32790 not n7914 ; n7914_not
g32791 not n1497 ; n1497_not
g32792 not n6258 ; n6258_not
g32793 not n9534 ; n9534_not
g32794 not n4872 ; n4872_not
g32795 not n7293 ; n7293_not
g32796 not n2775 ; n2775_not
g32797 not n3882 ; n3882_not
g32798 not n3936 ; n3936_not
g32799 not n3576 ; n3576_not
g32800 not n8535 ; n8535_not
g32801 not n9237 ; n9237_not
g32802 not n9813 ; n9813_not
g32803 not n3855 ; n3855_not
g32804 not n7158 ; n7158_not
g32805 not n9507 ; n9507_not
g32806 not n4188 ; n4188_not
g32807 not n8382 ; n8382_not
g32808 not n7950 ; n7950_not
g32809 not n4179 ; n4179_not
g32810 not n7167 ; n7167_not
g32811 not n2838 ; n2838_not
g32812 not n7149 ; n7149_not
g32813 not n6474 ; n6474_not
g32814 not n6087 ; n6087_not
g32815 not n7626 ; n7626_not
g32816 not n8391 ; n8391_not
g32817 not n8373 ; n8373_not
g32818 not n5466 ; n5466_not
g32819 not n9246 ; n9246_not
g32820 not n8544 ; n8544_not
g32821 not n7644 ; n7644_not
g32822 not n9192 ; n9192_not
g32823 not n3288 ; n3288_not
g32824 not n4269 ; n4269_not
g32825 not n5475 ; n5475_not
g32826 not n6096 ; n6096_not
g32827 not n4089 ; n4089_not
g32828 not n3873 ; n3873_not
g32829 not n8067 ; n8067_not
g32830 not n9282 ; n9282_not
g32831 not n9426 ; n9426_not
g32832 not n8517 ; n8517_not
g32833 not n8328 ; n8328_not
g32834 not n6069 ; n6069_not
g32835 not n9273 ; n9273_not
g32836 not n5628 ; n5628_not
g32837 not n1686 ; n1686_not
g32838 not n8508 ; n8508_not
g32839 not n2829 ; n2829_not
g32840 not n3567 ; n3567_not
g32841 not n5538 ; n5538_not
g32842 not n2739 ; n2739_not
g32843 not n5493 ; n5493_not
g32844 not n7176 ; n7176_not
g32845 not n4881 ; n4881_not
g32846 not n7185 ; n7185_not
g32847 not n3864 ; n3864_not
g32848 not n2694 ; n2694_not
g32849 not n7941 ; n7941_not
g32850 not n4098 ; n4098_not
g32851 not n1578 ; n1578_not
g32852 not n5394 ; n5394_not
g32853 not n7194 ; n7194_not
g32854 not n7383 ; n7383_not
g32855 not n6429 ; n6429_not
g32856 not n8526 ; n8526_not
g32857 not n6078 ; n6078_not
g32858 not n4854 ; n4854_not
g32859 not n6537 ; n6537_not
g32860 not n7554 ; n7554_not
g32861 not n6573 ; n6573_not
g32862 not n8751 ; n8751_not
g32863 not n1965 ; n1965_not
g32864 not n3396 ; n3396_not
g32865 not n9048 ; n9048_not
g32866 not n6294 ; n6294_not
g32867 not n4665 ; n4665_not
g32868 not n6744 ; n6744_not
g32869 not n2964 ; n2964_not
g32870 not n5952 ; n5952_not
g32871 not n4674 ; n4674_not
g32872 not n9183 ; n9183_not
g32873 not n2199 ; n2199_not
g32874 not n2973 ; n2973_not
g32875 not n9075 ; n9075_not
g32876 not n9363 ; n9363_not
g32877 not n9084 ; n9084_not
g32878 not n9372 ; n9372_not
g32879 not n6375 ; n6375_not
g32880 not n3387 ; n3387_not
g32881 not n6582 ; n6582_not
g32882 not n6717 ; n6717_not
g32883 not n3693 ; n3693_not
g32884 not n9066 ; n9066_not
g32885 not n9381 ; n9381_not
g32886 not n5655 ; n5655_not
g32887 not n4683 ; n4683_not
g32888 not n4782 ; n4782_not
g32889 not n6726 ; n6726_not
g32890 not n9390 ; n9390_not
g32891 not n2379 ; n2379_not
g32892 not n1299 ; n1299_not
g32893 not n6267 ; n6267_not
g32894 not n2388 ; n2388_not
g32895 not n8238 ; n8238_not
g32896 not n2397 ; n2397_not
g32897 not n7581 ; n7581_not
g32898 not n8148 ; n8148_not
g32899 not n1659 ; n1659_not
g32900 not n2946 ; n2946_not
g32901 not n7680 ; n7680_not
g32902 not n7743 ; n7743_not
g32903 not n8247 ; n8247_not
g32904 not n8940 ; n8940_not
g32905 not n6555 ; n6555_not
g32906 not n7572 ; n7572_not
g32907 not n8931 ; n8931_not
g32908 not n5088 ; n5088_not
g32909 not n6285 ; n6285_not
g32910 not n1677 ; n1677_not
g32911 not n8058 ; n8058_not
g32912 not n6753 ; n6753_not
g32913 not n9039 ; n9039_not
g32914 not n9408 ; n9408_not
g32915 not n1389 ; n1389_not
g32916 not n2289 ; n2289_not
g32917 not n7671 ; n7671_not
g32918 not n1668 ; n1668_not
g32919 not n6564 ; n6564_not
g32920 not n2298 ; n2298_not
g32921 not n7590 ; n7590_not
g32922 not n7806 ; n7806_not
g32923 not n6276 ; n6276_not
g32924 not n1947 ; n1947_not
g32925 not n4755 ; n4755_not
g32926 not n1695 ; n1695_not
g32927 not n7761 ; n7761_not
g32928 not n3378 ; n3378_not
g32929 not n8184 ; n8184_not
g32930 not n6636 ; n6636_not
g32931 not n4953 ; n4953_not
g32932 not n9624 ; n9624_not
g32933 not n6348 ; n6348_not
g32934 not n1956 ; n1956_not
g32935 not n7374 ; n7374_not
g32936 not n3675 ; n3675_not
g32937 not n4935 ; n4935_not
g32938 not n4737 ; n4737_not
g32939 not n4647 ; n4647_not
g32940 not n4773 ; n4773_not
g32941 not n8085 ; n8085_not
g32942 not n5916 ; n5916_not
g32943 not n6609 ; n6609_not
g32944 not n9336 ; n9336_not
g32945 not n4944 ; n4944_not
g32946 not n8094 ; n8094_not
g32947 not n1884 ; n1884_not
g32948 not n4764 ; n4764_not
g32949 not n6357 ; n6357_not
g32950 not n7653 ; n7653_not
g32951 not n6618 ; n6618_not
g32952 not n9147 ; n9147_not
g32953 not n1749 ; n1749_not
g32954 not n6627 ; n6627_not
g32955 not n9156 ; n9156_not
g32956 not n1938 ; n1938_not
g32957 not n9318 ; n9318_not
g32958 not n9057 ; n9057_not
g32959 not n9354 ; n9354_not
g32960 not n5745 ; n5745_not
g32961 not n6681 ; n6681_not
g32962 not n2991 ; n2991_not
g32963 not n9165 ; n9165_not
g32964 not n1992 ; n1992_not
g32965 not n3684 ; n3684_not
g32966 not n4971 ; n4971_not
g32967 not n9093 ; n9093_not
g32968 not n7617 ; n7617_not
g32969 not n5907 ; n5907_not
g32970 not n9633 ; n9633_not
g32971 not n8076 ; n8076_not
g32972 not n8166 ; n8166_not
g32973 not n5619 ; n5619_not
g32974 not n5637 ; n5637_not
g32975 not n9327 ; n9327_not
g32976 not n3369 ; n3369_not
g32977 not n4728 ; n4728_not
g32978 not n6654 ; n6654_not
g32979 not n9345 ; n9345_not
g32980 not n6591 ; n6591_not
g32981 not n7635 ; n7635_not
g32982 not n7770 ; n7770_not
g32983 not n6663 ; n6663_not
g32984 not n1974 ; n1974_not
g32985 not n6339 ; n6339_not
g32986 not n6672 ; n6672_not
g32987 not n4962 ; n4962_not
g32988 not n1983 ; n1983_not
g32989 not n7662 ; n7662_not
g32990 not n8139 ; n8139_not
g32991 not n8823 ; n8823_not
g32992 not n2469 ; n2469_not
g32993 not n5178 ; n5178_not
g32994 not n8805 ; n8805_not
g32995 not n8814 ; n8814_not
g32996 not n3459 ; n3459_not
g32997 not n5691 ; n5691_not
g32998 not n5169 ; n5169_not
g32999 not n5187 ; n5187_not
g33000 not n2487 ; n2487_not
g33001 not n9930 ; n9930_not
g33002 not n3639 ; n3639_not
g33003 not n3729 ; n3729_not
g33004 not n6852 ; n6852_not
g33005 not n8850 ; n8850_not
g33006 not n8661 ; n8661_not
g33007 not n6861 ; n6861_not
g33008 not n8841 ; n8841_not
g33009 not n6393 ; n6393_not
g33010 not n6870 ; n6870_not
g33011 not n7545 ; n7545_not
g33012 not n8832 ; n8832_not
g33013 not n7815 ; n7815_not
g33014 not n3585 ; n3585_not
g33015 not n8274 ; n8274_not
g33016 not n2919 ; n2919_not
g33017 not n4818 ; n4818_not
g33018 not n5970 ; n5970_not
g33019 not n8742 ; n8742_not
g33020 not n3297 ; n3297_not
g33021 not n9912 ; n9912_not
g33022 not n4746 ; n4746_not
g33023 not n8724 ; n8724_not
g33024 not n6519 ; n6519_not
g33025 not n4593 ; n4593_not
g33026 not n3747 ; n3747_not
g33027 not n3099 ; n3099_not
g33028 not n9921 ; n9921_not
g33029 not n4809 ; n4809_not
g33030 not n7527 ; n7527_not
g33031 not n5196 ; n5196_not
g33032 not n9903 ; n9903_not
g33033 not n8760 ; n8760_not
g33034 not n3756 ; n3756_not
g33035 not n9615 ; n9615_not
g33036 not n4584 ; n4584_not
g33037 not n6924 ; n6924_not
g33038 not n7518 ; n7518_not
g33039 not n1875 ; n1875_not
g33040 not n8049 ; n8049_not
g33041 not n5664 ; n5664_not
g33042 not n7563 ; n7563_not
g33043 not n4926 ; n4926_not
g33044 not n1893 ; n1893_not
g33045 not n5781 ; n5781_not
g33046 not n9723 ; n9723_not
g33047 not n9417 ; n9417_not
g33048 not n5943 ; n5943_not
g33049 not n5097 ; n5097_not
g33050 not n6834 ; n6834_not
g33051 not n5880 ; n5880_not
g33052 not n8256 ; n8256_not
g33053 not n6249 ; n6249_not
g33054 not n6816 ; n6816_not
g33055 not n9714 ; n9714_not
g33056 not n6546 ; n6546_not
g33057 not n4656 ; n4656_not
g33058 not n2928 ; n2928_not
g33059 not n5961 ; n5961_not
g33060 not n3594 ; n3594_not
g33061 not n5718 ; n5718_not
g33062 not n3379 ; n3379_not
g33063 not n3676 ; n3676_not
g33064 not n8419 ; n8419_not
g33065 not n7681 ; n7681_not
g33066 not n3757 ; n3757_not
g33067 not n5755 ; n5755_not
g33068 not n7834 ; n7834_not
g33069 not n3289 ; n3289_not
g33070 not n7807 ; n7807_not
g33071 not n8239 ; n8239_not
g33072 not n5728 ; n5728_not
g33073 not n2875 ; n2875_not
g33074 not n3586 ; n3586_not
g33075 not n8086 ; n8086_not
g33076 not n7465 ; n7465_not
g33077 not n8149 ; n8149_not
g33078 not n7528 ; n7528_not
g33079 not n9904 ; n9904_not
g33080 not n7924 ; n7924_not
g33081 not n9841 ; n9841_not
g33082 not n2794 ; n2794_not
g33083 not n5683 ; n5683_not
g33084 not n7438 ; n7438_not
g33085 not n7636 ; n7636_not
g33086 not n8176 ; n8176_not
g33087 not n7357 ; n7357_not
g33088 not n5656 ; n5656_not
g33089 not n7483 ; n7483_not
g33090 not n7627 ; n7627_not
g33091 not n7717 ; n7717_not
g33092 not n8293 ; n8293_not
g33093 not n8248 ; n8248_not
g33094 not n3883 ; n3883_not
g33095 not n8275 ; n8275_not
g33096 not n5791 ; n5791_not
g33097 not n7573 ; n7573_not
g33098 not n7654 ; n7654_not
g33099 not n5638 ; n5638_not
g33100 not n7339 ; n7339_not
g33101 not n7870 ; n7870_not
g33102 not n2938 ; n2938_not
g33103 not n7762 ; n7762_not
g33104 not n8284 ; n8284_not
g33105 not n3766 ; n3766_not
g33106 not n9913 ; n9913_not
g33107 not n5737 ; n5737_not
g33108 not n3775 ; n3775_not
g33109 not n7906 ; n7906_not
g33110 not n2992 ; n2992_not
g33111 not n8095 ; n8095_not
g33112 not n5764 ; n5764_not
g33113 not n7852 ; n7852_not
g33114 not n3874 ; n3874_not
g33115 not n3694 ; n3694_not
g33116 not n7348 ; n7348_not
g33117 not n8185 ; n8185_not
g33118 not n7168 ; n7168_not
g33119 not n9940 ; n9940_not
g33120 not n7915 ; n7915_not
g33121 not n2929 ; n2929_not
g33122 not n9814 ; n9814_not
g33123 not n3469 ; n3469_not
g33124 not n7645 ; n7645_not
g33125 not n7519 ; n7519_not
g33126 not n7492 ; n7492_not
g33127 not n8194 ; n8194_not
g33128 not n7825 ; n7825_not
g33129 not n9922 ; n9922_not
g33130 not n8167 ; n8167_not
g33131 not n7456 ; n7456_not
g33132 not n5773 ; n5773_not
g33133 not n3199 ; n3199_not
g33134 not n2848 ; n2848_not
g33135 not n7447 ; n7447_not
g33136 not n7267 ; n7267_not
g33137 not n3793 ; n3793_not
g33138 not n7582 ; n7582_not
g33139 not n8266 ; n8266_not
g33140 not n7546 ; n7546_not
g33141 not n7285 ; n7285_not
g33142 not n7942 ; n7942_not
g33143 not n7672 ; n7672_not
g33144 not n2974 ; n2974_not
g33145 not n7384 ; n7384_not
g33146 not n8068 ; n8068_not
g33147 not n3559 ; n3559_not
g33148 not n7816 ; n7816_not
g33149 not n3388 ; n3388_not
g33150 not n8374 ; n8374_not
g33151 not n9850 ; n9850_not
g33152 not n8257 ; n8257_not
g33153 not n5782 ; n5782_not
g33154 not n2857 ; n2857_not
g33155 not n3658 ; n3658_not
g33156 not n8356 ; n8356_not
g33157 not n7960 ; n7960_not
g33158 not n3487 ; n3487_not
g33159 not n2776 ; n2776_not
g33160 not n7951 ; n7951_not
g33161 not n7771 ; n7771_not
g33162 not n8383 ; n8383_not
g33163 not n8158 ; n8158_not
g33164 not n8365 ; n8365_not
g33165 not n9931 ; n9931_not
g33166 not n2965 ; n2965_not
g33167 not n7618 ; n7618_not
g33168 not n9643 ; n9643_not
g33169 not n7177 ; n7177_not
g33170 not n7663 ; n7663_not
g33171 not n2947 ; n2947_not
g33172 not n3739 ; n3739_not
g33173 not n7861 ; n7861_not
g33174 not n7708 ; n7708_not
g33175 not n3748 ; n3748_not
g33176 not n8329 ; n8329_not
g33177 not n7366 ; n7366_not
g33178 not n7474 ; n7474_not
g33179 not n5746 ; n5746_not
g33180 not n3568 ; n3568_not
g33181 not n7735 ; n7735_not
g33182 not n7690 ; n7690_not
g33183 not n7564 ; n7564_not
g33184 not n7780 ; n7780_not
g33185 not n3865 ; n3865_not
g33186 not n7609 ; n7609_not
g33187 not n2839 ; n2839_not
g33188 not n7375 ; n7375_not
g33189 not n3649 ; n3649_not
g33190 not n7591 ; n7591_not
g33191 not n7744 ; n7744_not
g33192 not n7537 ; n7537_not
g33193 not n8347 ; n8347_not
g33194 not n5809 ; n5809_not
g33195 not n3478 ; n3478_not
g33196 not n3856 ; n3856_not
g33197 not n8077 ; n8077_not
g33198 not n8338 ; n8338_not
g33199 not n5926 ; n5926_not
g33200 not n4819 ; n4819_not
g33201 not n6529 ; n6529_not
g33202 not n4747 ; n4747_not
g33203 not n1876 ; n1876_not
g33204 not n6259 ; n6259_not
g33205 not n6538 ; n6538_not
g33206 not n6547 ; n6547_not
g33207 not n4792 ; n4792_not
g33208 not n6556 ; n6556_not
g33209 not n1894 ; n1894_not
g33210 not n9193 ; n9193_not
g33211 not n6358 ; n6358_not
g33212 not n6349 ; n6349_not
g33213 not n9184 ; n9184_not
g33214 not n6628 ; n6628_not
g33215 not n6619 ; n6619_not
g33216 not n9652 ; n9652_not
g33217 not n9148 ; n9148_not
g33218 not n6574 ; n6574_not
g33219 not n4774 ; n4774_not
g33220 not n1939 ; n1939_not
g33221 not n4765 ; n4765_not
g33222 not n1885 ; n1885_not
g33223 not n5647 ; n5647_not
g33224 not n6592 ; n6592_not
g33225 not n9166 ; n9166_not
g33226 not n6583 ; n6583_not
g33227 not n4783 ; n4783_not
g33228 not n9175 ; n9175_not
g33229 not n9256 ; n9256_not
g33230 not n5935 ; n5935_not
g33231 not n9265 ; n9265_not
g33232 not n4864 ; n4864_not
g33233 not n6448 ; n6448_not
g33234 not n4873 ; n4873_not
g33235 not n1795 ; n1795_not
g33236 not n6439 ; n6439_not
g33237 not n9274 ; n9274_not
g33238 not n4882 ; n4882_not
g33239 not n9283 ; n9283_not
g33240 not n1786 ; n1786_not
g33241 not n4909 ; n4909_not
g33242 not n1867 ; n1867_not
g33243 not n4837 ; n4837_not
g33244 not n4828 ; n4828_not
g33245 not n9229 ; n9229_not
g33246 not n1858 ; n1858_not
g33247 not n1849 ; n1849_not
g33248 not n6493 ; n6493_not
g33249 not n9238 ; n9238_not
g33250 not n6484 ; n6484_not
g33251 not n4846 ; n4846_not
g33252 not n9247 ; n9247_not
g33253 not n6475 ; n6475_not
g33254 not n4855 ; n4855_not
g33255 not n5629 ; n5629_not
g33256 not n6466 ; n6466_not
g33257 not n6727 ; n6727_not
g33258 not n9058 ; n9058_not
g33259 not n9481 ; n9481_not
g33260 not n9670 ; n9670_not
g33261 not n4675 ; n4675_not
g33262 not n6745 ; n6745_not
g33263 not n6754 ; n6754_not
g33264 not n4666 ; n4666_not
g33265 not n6763 ; n6763_not
g33266 not n2299 ; n2299_not
g33267 not n9706 ; n9706_not
g33268 not n6772 ; n6772_not
g33269 not n2389 ; n2389_not
g33270 not n6844 ; n6844_not
g33271 not n9724 ; n9724_not
g33272 not n6835 ; n6835_not
g33273 not n5881 ; n5881_not
g33274 not n8914 ; n8914_not
g33275 not n6817 ; n6817_not
g33276 not n9715 ; n9715_not
g33277 not n4648 ; n4648_not
g33278 not n8932 ; n8932_not
g33279 not n2398 ; n2398_not
g33280 not n8950 ; n8950_not
g33281 not n8635 ; n8635_not
g33282 not n6790 ; n6790_not
g33283 not n8860 ; n8860_not
g33284 not n8851 ; n8851_not
g33285 not n6673 ; n6673_not
g33286 not n1975 ; n1975_not
g33287 not n6664 ; n6664_not
g33288 not n6376 ; n6376_not
g33289 not n4729 ; n4729_not
g33290 not n1966 ; n1966_not
g33291 not n6655 ; n6655_not
g33292 not n5719 ; n5719_not
g33293 not n6646 ; n6646_not
g33294 not n4738 ; n4738_not
g33295 not n9661 ; n9661_not
g33296 not n6637 ; n6637_not
g33297 not n4576 ; n4576_not
g33298 not n1948 ; n1948_not
g33299 not n4756 ; n4756_not
g33300 not n9067 ; n9067_not
g33301 not n6718 ; n6718_not
g33302 not n4693 ; n4693_not
g33303 not n9076 ; n9076_not
g33304 not n9085 ; n9085_not
g33305 not n4684 ; n4684_not
g33306 not n9094 ; n9094_not
g33307 not n6691 ; n6691_not
g33308 not n1993 ; n1993_not
g33309 not n5908 ; n5908_not
g33310 not n6682 ; n6682_not
g33311 not n6394 ; n6394_not
g33312 not n9472 ; n9472_not
g33313 not n5395 ; n5395_not
g33314 not n5980 ; n5980_not
g33315 not n5377 ; n5377_not
g33316 not n9463 ; n9463_not
g33317 not n5386 ; n5386_not
g33318 not n5098 ; n5098_not
g33319 not n9454 ; n9454_not
g33320 not n5368 ; n5368_not
g33321 not n9607 ; n9607_not
g33322 not n5359 ; n5359_not
g33323 not n1489 ; n1489_not
g33324 not n5962 ; n5962_not
g33325 not n9427 ; n9427_not
g33326 not n5692 ; n5692_not
g33327 not n9436 ; n9436_not
g33328 not n6196 ; n6196_not
g33329 not n6187 ; n6187_not
g33330 not n5971 ; n5971_not
g33331 not n5269 ; n5269_not
g33332 not n5278 ; n5278_not
g33333 not n6178 ; n6178_not
g33334 not n5287 ; n5287_not
g33335 not n6169 ; n6169_not
g33336 not n9445 ; n9445_not
g33337 not n5296 ; n5296_not
g33338 not n1588 ; n1588_not
g33339 not n9571 ; n9571_not
g33340 not n5539 ; n5539_not
g33341 not n5548 ; n5548_not
g33342 not n9517 ; n9517_not
g33343 not n5557 ; n5557_not
g33344 not n9562 ; n9562_not
g33345 not n5566 ; n5566_not
g33346 not n9553 ; n9553_not
g33347 not n5575 ; n5575_not
g33348 not n5485 ; n5485_not
g33349 not n9535 ; n9535_not
g33350 not n5584 ; n5584_not
g33351 not n1498 ; n1498_not
g33352 not n5593 ; n5593_not
g33353 not n5449 ; n5449_not
g33354 not n9490 ; n9490_not
g33355 not n5467 ; n5467_not
g33356 not n6097 ; n6097_not
g33357 not n9580 ; n9580_not
g33358 not n1579 ; n1579_not
g33359 not n9508 ; n9508_not
g33360 not n6088 ; n6088_not
g33361 not n5494 ; n5494_not
g33362 not n6079 ; n6079_not
g33363 not n4972 ; n4972_not
g33364 not n9355 ; n9355_not
g33365 not n9616 ; n9616_not
g33366 not n9346 ; n9346_not
g33367 not n6295 ; n6295_not
g33368 not n4945 ; n4945_not
g33369 not n9337 ; n9337_not
g33370 not n6367 ; n6367_not
g33371 not n1399 ; n1399_not
g33372 not n4918 ; n4918_not
g33373 not n1777 ; n1777_not
g33374 not n1768 ; n1768_not
g33375 not n9319 ; n9319_not
g33376 not n6385 ; n6385_not
g33377 not n4927 ; n4927_not
g33378 not n1759 ; n1759_not
g33379 not n9634 ; n9634_not
g33380 not n4936 ; n4936_not
g33381 not n9328 ; n9328_not
g33382 not n5944 ; n5944_not
g33383 not n1669 ; n1669_not
g33384 not n9625 ; n9625_not
g33385 not n5089 ; n5089_not
g33386 not n4963 ; n4963_not
g33387 not n9418 ; n9418_not
g33388 not n9409 ; n9409_not
g33389 not n9292 ; n9292_not
g33390 not n5179 ; n5179_not
g33391 not n5188 ; n5188_not
g33392 not n5953 ; n5953_not
g33393 not n9364 ; n9364_not
g33394 not n9373 ; n9373_not
g33395 not n4990 ; n4990_not
g33396 not n1687 ; n1687_not
g33397 not n9391 ; n9391_not
g33398 not n1678 ; n1678_not
g33399 not n6286 ; n6286_not
g33400 not n6277 ; n6277_not
g33401 not n6268 ; n6268_not
g33402 not n6862 ; n6862_not
g33403 not n8653 ; n8653_not
g33404 not n8527 ; n8527_not
g33405 not n8509 ; n8509_not
g33406 not n8644 ; n8644_not
g33407 not n7186 ; n7186_not
g33408 not n5458 ; n5458_not
g33409 not n2596 ; n2596_not
g33410 not n4099 ; n4099_not
g33411 not n8626 ; n8626_not
g33412 not n9742 ; n9742_not
g33413 not n9751 ; n9751_not
g33414 not n3955 ; n3955_not
g33415 not n5863 ; n5863_not
g33416 not n7249 ; n7249_not
g33417 not n9733 ; n9733_not
g33418 not n3973 ; n3973_not
g33419 not n6952 ; n6952_not
g33420 not n8716 ; n8716_not
g33421 not n8491 ; n8491_not
g33422 not n2569 ; n2569_not
g33423 not n5818 ; n5818_not
g33424 not n2749 ; n2749_not
g33425 not n8707 ; n8707_not
g33426 not n3991 ; n3991_not
g33427 not n3982 ; n3982_not
g33428 not n6961 ; n6961_not
g33429 not n2578 ; n2578_not
g33430 not n2668 ; n2668_not
g33431 not n3937 ; n3937_not
g33432 not n8482 ; n8482_not
g33433 not n3928 ; n3928_not
g33434 not n8518 ; n8518_not
g33435 not n8671 ; n8671_not
g33436 not n2695 ; n2695_not
g33437 not n5854 ; n5854_not
g33438 not n8581 ; n8581_not
g33439 not n7069 ; n7069_not
g33440 not n9805 ; n9805_not
g33441 not n4288 ; n4288_not
g33442 not n2677 ; n2677_not
g33443 not n4297 ; n4297_not
g33444 not n4396 ; n4396_not
g33445 not n7078 ; n7078_not
g33446 not n8572 ; n8572_not
g33447 not n8554 ; n8554_not
g33448 not n4387 ; n4387_not
g33449 not n5845 ; n5845_not
g33450 not n8563 ; n8563_not
g33451 not n7096 ; n7096_not
g33452 not n4369 ; n4369_not
g33453 not n4378 ; n4378_not
g33454 not n4567 ; n4567_not
g33455 not n4558 ; n4558_not
g33456 not n6826 ; n6826_not
g33457 not n5665 ; n5665_not
g33458 not n9760 ; n9760_not
g33459 not n5836 ; n5836_not
g33460 not n7159 ; n7159_not
g33461 not n8608 ; n8608_not
g33462 not n2659 ; n2659_not
g33463 not n4189 ; n4189_not
g33464 not n2686 ; n2686_not
g33465 not n9382 ; n9382_not
g33466 not n6934 ; n6934_not
g33467 not n5674 ; n5674_not
g33468 not n4486 ; n4486_not
g33469 not n8545 ; n8545_not
g33470 not n4279 ; n4279_not
g33471 not n4477 ; n4477_not
g33472 not n8590 ; n8590_not
g33473 not n4468 ; n4468_not
g33474 not n8833 ; n8833_not
g33475 not n8815 ; n8815_not
g33476 not n8446 ; n8446_not
g33477 not n2479 ; n2479_not
g33478 not n8806 ; n8806_not
g33479 not n2488 ; n2488_not
g33480 not n3946 ; n3946_not
g33481 not n6907 ; n6907_not
g33482 not n8770 ; n8770_not
g33483 not n2767 ; n2767_not
g33484 not n8761 ; n8761_not
g33485 not n7276 ; n7276_not
g33486 not n2758 ; n2758_not
g33487 not n2785 ; n2785_not
g33488 not n8428 ; n8428_not
g33489 not n8905 ; n8905_not
g33490 not n3892 ; n3892_not
g33491 not n6853 ; n6853_not
g33492 not n8662 ; n8662_not
g33493 not n3838 ; n3838_not
g33494 not n9823 ; n9823_not
g33495 not n8842 ; n8842_not
g33496 not n8824 ; n8824_not
g33497 not n3919 ; n3919_not
g33498 not n7087 ; n7087_not
g33499 not n7294 ; n7294_not
g33500 not n6871 ; n6871_not
g33501 not n8464 ; n8464_not
g33502 not n8752 ; n8752_not
g33503 not n6916 ; n6916_not
g33504 not n4585 ; n4585_not
g33505 not n6925 ; n6925_not
g33506 not n3964 ; n3964_not
g33507 not n8743 ; n8743_not
g33508 not n8473 ; n8473_not
g33509 not n7258 ; n7258_not
g33510 not n8734 ; n8734_not
g33511 not n8725 ; n8725_not
g33512 not n6943 ; n6943_not
g33513 not n9527 ; n9527_not
g33514 not n3488 ; n3488_not
g33515 not n9428 ; n9428_not
g33516 not n9365 ; n9365_not
g33517 not n3299 ; n3299_not
g33518 not n3389 ; n3389_not
g33519 not n9860 ; n9860_not
g33520 not n8492 ; n8492_not
g33521 not n8528 ; n8528_not
g33522 not n2795 ; n2795_not
g33523 not n9518 ; n9518_not
g33524 not n8069 ; n8069_not
g33525 not n9383 ; n9383_not
g33526 not n2759 ; n2759_not
g33527 not n2678 ; n2678_not
g33528 not n9608 ; n9608_not
g33529 not n9392 ; n9392_not
g33530 not n8546 ; n8546_not
g33531 not n9437 ; n9437_not
g33532 not n8483 ; n8483_not
g33533 not n9536 ; n9536_not
g33534 not n9356 ; n9356_not
g33535 not n7907 ; n7907_not
g33536 not n7709 ; n7709_not
g33537 not n3578 ; n3578_not
g33538 not n9455 ; n9455_not
g33539 not n1499 ; n1499_not
g33540 not n2786 ; n2786_not
g33541 not n8429 ; n8429_not
g33542 not n9824 ; n9824_not
g33543 not n7745 ; n7745_not
g33544 not n9464 ; n9464_not
g33545 not n2777 ; n2777_not
g33546 not n8438 ; n8438_not
g33547 not n9554 ; n9554_not
g33548 not n7916 ; n7916_not
g33549 not n9374 ; n9374_not
g33550 not n2687 ; n2687_not
g33551 not n9509 ; n9509_not
g33552 not n8465 ; n8465_not
g33553 not n9590 ; n9590_not
g33554 not n7943 ; n7943_not
g33555 not n9617 ; n9617_not
g33556 not n9842 ; n9842_not
g33557 not n9572 ; n9572_not
g33558 not n1589 ; n1589_not
g33559 not n7961 ; n7961_not
g33560 not n7844 ; n7844_not
g33561 not n9419 ; n9419_not
g33562 not n8384 ; n8384_not
g33563 not n8519 ; n8519_not
g33564 not n9581 ; n9581_not
g33565 not n2696 ; n2696_not
g33566 not n9680 ; n9680_not
g33567 not n8447 ; n8447_not
g33568 not n9473 ; n9473_not
g33569 not n1679 ; n1679_not
g33570 not n3398 ; n3398_not
g33571 not n8375 ; n8375_not
g33572 not n9851 ; n9851_not
g33573 not n8537 ; n8537_not
g33574 not n7970 ; n7970_not
g33575 not n9491 ; n9491_not
g33576 not n9815 ; n9815_not
g33577 not n9626 ; n9626_not
g33578 not n9446 ; n9446_not
g33579 not n8339 ; n8339_not
g33580 not n3479 ; n3479_not
g33581 not n7934 ; n7934_not
g33582 not n7952 ; n7952_not
g33583 not n1985 ; n1985_not
g33584 not n2498 ; n2498_not
g33585 not n8753 ; n8753_not
g33586 not n1994 ; n1994_not
g33587 not n8195 ; n8195_not
g33588 not n2984 ; n2984_not
g33589 not n9095 ; n9095_not
g33590 not n8762 ; n8762_not
g33591 not n8744 ; n8744_not
g33592 not n9068 ; n9068_not
g33593 not n9086 ; n9086_not
g33594 not n2975 ; n2975_not
g33595 not n8780 ; n8780_not
g33596 not n9077 ; n9077_not
g33597 not n2489 ; n2489_not
g33598 not n9923 ; n9923_not
g33599 not n8708 ; n8708_not
g33600 not n9149 ; n9149_not
g33601 not n9734 ; n9734_not
g33602 not n8285 ; n8285_not
g33603 not n9653 ; n9653_not
g33604 not n8717 ; n8717_not
g33605 not n1949 ; n1949_not
g33606 not n9338 ; n9338_not
g33607 not n9662 ; n9662_not
g33608 not n8186 ; n8186_not
g33609 not n8726 ; n8726_not
g33610 not n8735 ; n8735_not
g33611 not n2993 ; n2993_not
g33612 not n1967 ; n1967_not
g33613 not n8276 ; n8276_not
g33614 not n9914 ; n9914_not
g33615 not n8843 ; n8843_not
g33616 not n8951 ; n8951_not
g33617 not n8249 ; n8249_not
g33618 not n8933 ; n8933_not
g33619 not n2939 ; n2939_not
g33620 not n8852 ; n8852_not
g33621 not n8924 ; n8924_not
g33622 not n2399 ; n2399_not
g33623 not n9932 ; n9932_not
g33624 not n8915 ; n8915_not
g33625 not n8870 ; n8870_not
g33626 not n8258 ; n8258_not
g33627 not n8573 ; n8573_not
g33628 not n8906 ; n8906_not
g33629 not n9941 ; n9941_not
g33630 not n8807 ; n8807_not
g33631 not n9950 ; n9950_not
g33632 not n9059 ; n9059_not
g33633 not n2849 ; n2849_not
g33634 not n2966 ; n2966_not
g33635 not n8816 ; n8816_not
g33636 not n9725 ; n9725_not
g33637 not n2957 ; n2957_not
g33638 not n8825 ; n8825_not
g33639 not n9707 ; n9707_not
g33640 not n2948 ; n2948_not
g33641 not n8834 ; n8834_not
g33642 not n8267 ; n8267_not
g33643 not n8960 ; n8960_not
g33644 not n9716 ; n9716_not
g33645 not n2858 ; n2858_not
g33646 not n1787 ; n1787_not
g33647 not n9293 ; n9293_not
g33648 not n2669 ; n2669_not
g33649 not n9275 ; n9275_not
g33650 not n9284 ; n9284_not
g33651 not n9770 ; n9770_not
g33652 not n9761 ; n9761_not
g33653 not n1796 ; n1796_not
g33654 not n9905 ; n9905_not
g33655 not n8348 ; n8348_not
g33656 not n9257 ; n9257_not
g33657 not n8609 ; n8609_not
g33658 not n9248 ; n9248_not
g33659 not n9329 ; n9329_not
g33660 not n1697 ; n1697_not
g33661 not n9347 ; n9347_not
g33662 not n8087 ; n8087_not
g33663 not n8564 ; n8564_not
g33664 not n8096 ; n8096_not
g33665 not n8078 ; n8078_not
g33666 not n8582 ; n8582_not
g33667 not n8366 ; n8366_not
g33668 not n9635 ; n9635_not
g33669 not n1769 ; n1769_not
g33670 not n1778 ; n1778_not
g33671 not n8591 ; n8591_not
g33672 not n8663 ; n8663_not
g33673 not n2876 ; n2876_not
g33674 not n9185 ; n9185_not
g33675 not n2894 ; n2894_not
g33676 not n8672 ; n8672_not
g33677 not n8159 ; n8159_not
g33678 not n9176 ; n9176_not
g33679 not n2579 ; n2579_not
g33680 not n9167 ; n9167_not
g33681 not n8690 ; n8690_not
g33682 not n8294 ; n8294_not
g33683 not n8168 ; n8168_not
g33684 not n8177 ; n8177_not
g33685 not n2867 ; n2867_not
g33686 not n9752 ; n9752_not
g33687 not n9239 ; n9239_not
g33688 not n9743 ; n9743_not
g33689 not n9644 ; n9644_not
g33690 not n1859 ; n1859_not
g33691 not n8627 ; n8627_not
g33692 not n1868 ; n1868_not
g33693 not n2597 ; n2597_not
g33694 not n8636 ; n8636_not
g33695 not n1886 ; n1886_not
g33696 not n8645 ; n8645_not
g33697 not n2588 ; n2588_not
g33698 not n2885 ; n2885_not
g33699 not n1895 ; n1895_not
g33700 not n6962 ; n6962_not
g33701 not n5369 ; n5369_not
g33702 not n4298 ; n4298_not
g33703 not n6395 ; n6395_not
g33704 not n4649 ; n4649_not
g33705 not n3875 ; n3875_not
g33706 not n4379 ; n4379_not
g33707 not n6809 ; n6809_not
g33708 not n7754 ; n7754_not
g33709 not n5594 ; n5594_not
g33710 not n7097 ; n7097_not
g33711 not n6791 ; n6791_not
g33712 not n6674 ; n6674_not
g33713 not n4388 ; n4388_not
g33714 not n7547 ; n7547_not
g33715 not n7763 ; n7763_not
g33716 not n7259 ; n7259_not
g33717 not n7673 ; n7673_not
g33718 not n5783 ; n5783_not
g33719 not n5459 ; n5459_not
g33720 not n6692 ; n6692_not
g33721 not n6872 ; n6872_not
g33722 not n3893 ; n3893_not
g33723 not n3668 ; n3668_not
g33724 not n3659 ; n3659_not
g33725 not n7664 ; n7664_not
g33726 not n7718 ; n7718_not
g33727 not n6773 ; n6773_not
g33728 not n5648 ; n5648_not
g33729 not n6881 ; n6881_not
g33730 not n6746 ; n6746_not
g33731 not n6683 ; n6683_not
g33732 not n4883 ; n4883_not
g33733 not n7565 ; n7565_not
g33734 not n7556 ; n7556_not
g33735 not n7736 ; n7736_not
g33736 not n3767 ; n3767_not
g33737 not n5738 ; n5738_not
g33738 not n4748 ; n4748_not
g33739 not n6629 ; n6629_not
g33740 not n4757 ; n4757_not
g33741 not n4469 ; n4469_not
g33742 not n5774 ; n5774_not
g33743 not n5297 ; n5297_not
g33744 not n7358 ; n7358_not
g33745 not n3776 ; n3776_not
g33746 not n5288 ; n5288_not
g33747 not n4766 ; n4766_not
g33748 not n6908 ; n6908_not
g33749 not n7808 ; n7808_not
g33750 not n4487 ; n4487_not
g33751 not n3587 ; n3587_not
g33752 not n3884 ; n3884_not
g33753 not n6665 ; n6665_not
g33754 not n7079 ; n7079_not
g33755 not n7538 ; n7538_not
g33756 not n6890 ; n6890_not
g33757 not n3749 ; n3749_not
g33758 not n4397 ; n4397_not
g33759 not n5846 ; n5846_not
g33760 not n6656 ; n6656_not
g33761 not n7529 ; n7529_not
g33762 not n3758 ; n3758_not
g33763 not n7781 ; n7781_not
g33764 not n5675 ; n5675_not
g33765 not n6647 ; n6647_not
g33766 not n5558 ; n5558_not
g33767 not n7385 ; n7385_not
g33768 not n7628 ; n7628_not
g33769 not n7637 ; n7637_not
g33770 not n7277 ; n7277_not
g33771 not n6737 ; n6737_not
g33772 not n6845 ; n6845_not
g33773 not n5855 ; n5855_not
g33774 not n6971 ; n6971_not
g33775 not n6728 ; n6728_not
g33776 not n7655 ; n7655_not
g33777 not n7646 ; n7646_not
g33778 not n5396 ; n5396_not
g33779 not n6548 ; n6548_not
g33780 not n6764 ; n6764_not
g33781 not n3956 ; n3956_not
g33782 not n4676 ; n4676_not
g33783 not n4694 ; n4694_not
g33784 not n7619 ; n7619_not
g33785 not n5873 ; n5873_not
g33786 not n7268 ; n7268_not
g33787 not n5837 ; n5837_not
g33788 not n3695 ; n3695_not
g33789 not n6449 ; n6449_not
g33790 not n6755 ; n6755_not
g33791 not n3965 ; n3965_not
g33792 not n5189 ; n5189_not
g33793 not n5576 ; n5576_not
g33794 not n7088 ; n7088_not
g33795 not n4973 ; n4973_not
g33796 not n3938 ; n3938_not
g33797 not n3677 ; n3677_not
g33798 not n4658 ; n4658_not
g33799 not n5378 ; n5378_not
g33800 not n4991 ; n4991_not
g33801 not n7682 ; n7682_not
g33802 not n7196 ; n7196_not
g33803 not n6836 ; n6836_not
g33804 not n7178 ; n7178_not
g33805 not n5567 ; n5567_not
g33806 not n7295 ; n7295_not
g33807 not n7187 ; n7187_not
g33808 not n4667 ; n4667_not
g33809 not n7169 ; n7169_not
g33810 not n3929 ; n3929_not
g33811 not n4199 ; n4199_not
g33812 not n6827 ; n6827_not
g33813 not n4685 ; n4685_not
g33814 not n4919 ; n4919_not
g33815 not n7592 ; n7592_not
g33816 not n3983 ; n3983_not
g33817 not n6719 ; n6719_not
g33818 not n4982 ; n4982_not
g33819 not n3992 ; n3992_not
g33820 not n3947 ; n3947_not
g33821 not n7286 ; n7286_not
g33822 not n6854 ; n6854_not
g33823 not n7583 ; n7583_not
g33824 not n3794 ; n3794_not
g33825 not n5387 ; n5387_not
g33826 not n5666 ; n5666_not
g33827 not n5981 ; n5981_not
g33828 not n5909 ; n5909_not
g33829 not n6485 ; n6485_not
g33830 not n7871 ; n7871_not
g33831 not n6089 ; n6089_not
g33832 not n3848 ; n3848_not
g33833 not n6863 ; n6863_not
g33834 not n4838 ; n4838_not
g33835 not n6368 ; n6368_not
g33836 not n4865 ; n4865_not
g33837 not n3839 ; n3839_not
g33838 not n5963 ; n5963_not
g33839 not n4586 ; n4586_not
g33840 not n5756 ; n5756_not
g33841 not n6917 ; n6917_not
g33842 not n5927 ; n5927_not
g33843 not n5990 ; n5990_not
g33844 not n6980 ; n6980_not
g33845 not n4793 ; n4793_not
g33846 not n4928 ; n4928_not
g33847 not n3857 ; n3857_not
g33848 not n6539 ; n6539_not
g33849 not n7484 ; n7484_not
g33850 not n6458 ; n6458_not
g33851 not n5765 ; n5765_not
g33852 not n6467 ; n6467_not
g33853 not n5495 ; n5495_not
g33854 not n4829 ; n4829_not
g33855 not n7475 ; n7475_not
g33856 not n3785 ; n3785_not
g33857 not n6269 ; n6269_not
g33858 not n6278 ; n6278_not
g33859 not n6935 ; n6935_not
g33860 not n5729 ; n5729_not
g33861 not n6476 ; n6476_not
g33862 not n6638 ; n6638_not
g33863 not n4856 ; n4856_not
g33864 not n7457 ; n7457_not
g33865 not n6953 ; n6953_not
g33866 not n6287 ; n6287_not
g33867 not n6944 ; n6944_not
g33868 not n5486 ; n5486_not
g33869 not n5657 ; n5657_not
g33870 not n6926 ; n6926_not
g33871 not n5972 ; n5972_not
g33872 not n5549 ; n5549_not
g33873 not n7880 ; n7880_not
g33874 not n7439 ; n7439_not
g33875 not n4946 ; n4946_not
g33876 not n6494 ; n6494_not
g33877 not n4847 ; n4847_not
g33878 not n4964 ; n4964_not
g33879 not n6359 ; n6359_not
g33880 not n6179 ; n6179_not
g33881 not n7466 ; n7466_not
g33882 not n5792 ; n5792_not
g33883 not n4577 ; n4577_not
g33884 not n5279 ; n5279_not
g33885 not n7376 ; n7376_not
g33886 not n6584 ; n6584_not
g33887 not n6386 ; n6386_not
g33888 not n6575 ; n6575_not
g33889 not n3866 ; n3866_not
g33890 not n4874 ; n4874_not
g33891 not n7853 ; n7853_not
g33892 not n5864 ; n5864_not
g33893 not n4784 ; n4784_not
g33894 not n5693 ; n5693_not
g33895 not n5828 ; n5828_not
g33896 not n4775 ; n4775_not
g33897 not n7817 ; n7817_not
g33898 not n6098 ; n6098_not
g33899 not n5639 ; n5639_not
g33900 not n7772 ; n7772_not
g33901 not n6782 ; n6782_not
g33902 not n6593 ; n6593_not
g33903 not n7835 ; n7835_not
g33904 not n5468 ; n5468_not
g33905 not n7826 ; n7826_not
g33906 not n7349 ; n7349_not
g33907 not n5882 ; n5882_not
g33908 not n7367 ; n7367_not
g33909 not n6296 ; n6296_not
g33910 not n6197 ; n6197_not
g33911 not n5945 ; n5945_not
g33912 not n6557 ; n6557_not
g33913 not n7493 ; n7493_not
g33914 not n5684 ; n5684_not
g33915 not n7394 ; n7394_not
g33916 not n5954 ; n5954_not
g33917 not n6188 ; n6188_not
g33918 not n6377 ; n6377_not
g33919 not n5819 ; n5819_not
g33920 not n6846 ; n6846_not
g33921 not n4659 ; n4659_not
g33922 not n3858 ; n3858_not
g33923 not n2778 ; n2778_not
g33924 not n6792 ; n6792_not
g33925 not n6828 ; n6828_not
g33926 not n8385 ; n8385_not
g33927 not n2796 ; n2796_not
g33928 not n4947 ; n4947_not
g33929 not n8367 ; n8367_not
g33930 not n9348 ; n9348_not
g33931 not n3948 ; n3948_not
g33932 not n5955 ; n5955_not
g33933 not n5487 ; n5487_not
g33934 not n7395 ; n7395_not
g33935 not n7359 ; n7359_not
g33936 not n5928 ; n5928_not
g33937 not n8358 ; n8358_not
g33938 not n5478 ; n5478_not
g33939 not n1689 ; n1689_not
g33940 not n9483 ; n9483_not
g33941 not n8925 ; n8925_not
g33942 not n8943 ; n8943_not
g33943 not n3777 ; n3777_not
g33944 not n7269 ; n7269_not
g33945 not n3939 ; n3939_not
g33946 not n8934 ; n8934_not
g33947 not n8394 ; n8394_not
g33948 not n3885 ; n3885_not
g33949 not n4956 ; n4956_not
g33950 not n9771 ; n9771_not
g33951 not n4884 ; n4884_not
g33952 not n7296 ; n7296_not
g33953 not n3876 ; n3876_not
g33954 not n9492 ; n9492_not
g33955 not n6099 ; n6099_not
g33956 not n8448 ; n8448_not
g33957 not n8907 ; n8907_not
g33958 not n5469 ; n5469_not
g33959 not n7368 ; n7368_not
g33960 not n3894 ; n3894_not
g33961 not n5919 ; n5919_not
g33962 not n8457 ; n8457_not
g33963 not n8439 ; n8439_not
g33964 not n8952 ; n8952_not
g33965 not n3867 ; n3867_not
g33966 not n3849 ; n3849_not
g33967 not n7278 ; n7278_not
g33968 not n8376 ; n8376_not
g33969 not n7377 ; n7377_not
g33970 not n8628 ; n8628_not
g33971 not n6990 ; n6990_not
g33972 not n8781 ; n8781_not
g33973 not n6909 ; n6909_not
g33974 not n5982 ; n5982_not
g33975 not n9438 ; n9438_not
g33976 not n6189 ; n6189_not
g33977 not n6198 ; n6198_not
g33978 not n2589 ; n2589_not
g33979 not n9384 ; n9384_not
g33980 not n5685 ; n5685_not
g33981 not n8646 ; n8646_not
g33982 not n6981 ; n6981_not
g33983 not n8772 ; n8772_not
g33984 not n9843 ; n9843_not
g33985 not n9681 ; n9681_not
g33986 not n4488 ; n4488_not
g33987 not n5838 ; n5838_not
g33988 not n4497 ; n4497_not
g33989 not n5676 ; n5676_not
g33990 not n2598 ; n2598_not
g33991 not n5829 ; n5829_not
g33992 not n4389 ; n4389_not
g33993 not n6756 ; n6756_not
g33994 not n9816 ; n9816_not
g33995 not n6837 ; n6837_not
g33996 not n4578 ; n4578_not
g33997 not n6297 ; n6297_not
g33998 not n9852 ; n9852_not
g33999 not n9393 ; n9393_not
g34000 not n8619 ; n8619_not
g34001 not n1599 ; n1599_not
g34002 not n6918 ; n6918_not
g34003 not n6927 ; n6927_not
g34004 not n8691 ; n8691_not
g34005 not n4857 ; n4857_not
g34006 not n6963 ; n6963_not
g34007 not n2499 ; n2499_not
g34008 not n8745 ; n8745_not
g34009 not n9825 ; n9825_not
g34010 not n8709 ; n8709_not
g34011 not n6954 ; n6954_not
g34012 not n6279 ; n6279_not
g34013 not n8736 ; n8736_not
g34014 not n6936 ; n6936_not
g34015 not n9834 ; n9834_not
g34016 not n8727 ; n8727_not
g34017 not n7449 ; n7449_not
g34018 not n9429 ; n9429_not
g34019 not n6684 ; n6684_not
g34020 not n5199 ; n5199_not
g34021 not n8664 ; n8664_not
g34022 not n8754 ; n8754_not
g34023 not n5739 ; n5739_not
g34024 not n8763 ; n8763_not
g34025 not n6972 ; n6972_not
g34026 not n5694 ; n5694_not
g34027 not n4587 ; n4587_not
g34028 not n5649 ; n5649_not
g34029 not n9663 ; n9663_not
g34030 not n4938 ; n4938_not
g34031 not n8682 ; n8682_not
g34032 not n5856 ; n5856_not
g34033 not n3984 ; n3984_not
g34034 not n9096 ; n9096_not
g34035 not n8862 ; n8862_not
g34036 not n3993 ; n3993_not
g34037 not n4983 ; n4983_not
g34038 not n5388 ; n5388_not
g34039 not n9366 ; n9366_not
g34040 not n2679 ; n2679_not
g34041 not n8844 ; n8844_not
g34042 not n2697 ; n2697_not
g34043 not n7197 ; n7197_not
g34044 not n8673 ; n8673_not
g34045 not n8529 ; n8529_not
g34046 not n7188 ; n7188_not
g34047 not n7179 ; n7179_not
g34048 not n3975 ; n3975_not
g34049 not n9780 ; n9780_not
g34050 not n8169 ; n8169_not
g34051 not n8466 ; n8466_not
g34052 not n1698 ; n1698_not
g34053 not n4965 ; n4965_not
g34054 not n3966 ; n3966_not
g34055 not n3957 ; n3957_not
g34056 not n4974 ; n4974_not
g34057 not n8484 ; n8484_not
g34058 not n9465 ; n9465_not
g34059 not n9474 ; n9474_not
g34060 not n8493 ; n8493_not
g34061 not n5397 ; n5397_not
g34062 not n8871 ; n8871_not
g34063 not n8817 ; n8817_not
g34064 not n8259 ; n8259_not
g34065 not n5298 ; n5298_not
g34066 not n4398 ; n4398_not
g34067 not n9861 ; n9861_not
g34068 not n8583 ; n8583_not
g34069 not n8808 ; n8808_not
g34070 not n4596 ; n4596_not
g34071 not n9654 ; n9654_not
g34072 not n4479 ; n4479_not
g34073 not n8592 ; n8592_not
g34074 not n6594 ; n6594_not
g34075 not n5289 ; n5289_not
g34076 not n6774 ; n6774_not
g34077 not n5379 ; n5379_not
g34078 not n8538 ; n8538_not
g34079 not n9375 ; n9375_not
g34080 not n8835 ; n8835_not
g34081 not n6864 ; n6864_not
g34082 not n5847 ; n5847_not
g34083 not n6873 ; n6873_not
g34084 not n8547 ; n8547_not
g34085 not n9456 ; n9456_not
g34086 not n6882 ; n6882_not
g34087 not n8826 ; n8826_not
g34088 not n8556 ; n8556_not
g34089 not n4299 ; n4299_not
g34090 not n7098 ; n7098_not
g34091 not n7089 ; n7089_not
g34092 not n8565 ; n8565_not
g34093 not n9942 ; n9942_not
g34094 not n1959 ; n1959_not
g34095 not n7782 ; n7782_not
g34096 not n6648 ; n6648_not
g34097 not n5775 ; n5775_not
g34098 not n8079 ; n8079_not
g34099 not n7773 ; n7773_not
g34100 not n1968 ; n1968_not
g34101 not n8088 ; n8088_not
g34102 not n9555 ; n9555_not
g34103 not n9726 ; n9726_not
g34104 not n5595 ; n5595_not
g34105 not n7755 ; n7755_not
g34106 not n8097 ; n8097_not
g34107 not n6675 ; n6675_not
g34108 not n1986 ; n1986_not
g34109 not n9933 ; n9933_not
g34110 not n7548 ; n7548_not
g34111 not n4875 ; n4875_not
g34112 not n7917 ; n7917_not
g34113 not n7836 ; n7836_not
g34114 not n7827 ; n7827_not
g34115 not n4758 ; n4758_not
g34116 not n9159 ; n9159_not
g34117 not n4776 ; n4776_not
g34118 not n3588 ; n3588_not
g34119 not n7809 ; n7809_not
g34120 not n6585 ; n6585_not
g34121 not n3597 ; n3597_not
g34122 not n4767 ; n4767_not
g34123 not n9276 ; n9276_not
g34124 not n9951 ; n9951_not
g34125 not n3399 ; n3399_not
g34126 not n4749 ; n4749_not
g34127 not n6639 ; n6639_not
g34128 not n9087 ; n9087_not
g34129 not n9924 ; n9924_not
g34130 not n1788 ; n1788_not
g34131 not n7674 ; n7674_not
g34132 not n5874 ; n5874_not
g34133 not n4695 ; n4695_not
g34134 not n9078 ; n9078_not
g34135 not n9915 ; n9915_not
g34136 not n9168 ; n9168_not
g34137 not n9537 ; n9537_not
g34138 not n9069 ; n9069_not
g34139 not n3669 ; n3669_not
g34140 not n9294 ; n9294_not
g34141 not n7737 ; n7737_not
g34142 not n7575 ; n7575_not
g34143 not n7728 ; n7728_not
g34144 not n7719 ; n7719_not
g34145 not n5937 ; n5937_not
g34146 not n1995 ; n1995_not
g34147 not n7692 ; n7692_not
g34148 not n6693 ; n6693_not
g34149 not n5784 ; n5784_not
g34150 not n2967 ; n2967_not
g34151 not n1797 ; n1797_not
g34152 not n4893 ; n4893_not
g34153 not n7683 ; n7683_not
g34154 not n9546 ; n9546_not
g34155 not n6486 ; n6486_not
g34156 not n5964 ; n5964_not
g34157 not n5973 ; n5973_not
g34158 not n7935 ; n7935_not
g34159 not n9609 ; n9609_not
g34160 not n6477 ; n6477_not
g34161 not n6495 ; n6495_not
g34162 not n7944 ; n7944_not
g34163 not n7872 ; n7872_not
g34164 not n4839 ; n4839_not
g34165 not n7953 ; n7953_not
g34166 not n5757 ; n5757_not
g34167 not n7962 ; n7962_not
g34168 not n5892 ; n5892_not
g34169 not n3579 ; n3579_not
g34170 not n7908 ; n7908_not
g34171 not n7746 ; n7746_not
g34172 not n6468 ; n6468_not
g34173 not n9744 ; n9744_not
g34174 not n9762 ; n9762_not
g34175 not n9618 ; n9618_not
g34176 not n7890 ; n7890_not
g34177 not n9258 ; n9258_not
g34178 not n9249 ; n9249_not
g34179 not n4848 ; n4848_not
g34180 not n8916 ; n8916_not
g34181 not n7926 ; n7926_not
g34182 not n9708 ; n9708_not
g34183 not n9195 ; n9195_not
g34184 not n6558 ; n6558_not
g34185 not n9177 ; n9177_not
g34186 not n9186 ; n9186_not
g34187 not n6567 ; n6567_not
g34188 not n5991 ; n5991_not
g34189 not n7854 ; n7854_not
g34190 not n4785 ; n4785_not
g34191 not n6576 ; n6576_not
g34192 not n3498 ; n3498_not
g34193 not n1896 ; n1896_not
g34194 not n9717 ; n9717_not
g34195 not n3489 ; n3489_not
g34196 not n7845 ; n7845_not
g34197 not n5883 ; n5883_not
g34198 not n9627 ; n9627_not
g34199 not n6459 ; n6459_not
g34200 not n1869 ; n1869_not
g34201 not n4866 ; n4866_not
g34202 not n1887 ; n1887_not
g34203 not n9960 ; n9960_not
g34204 not n7980 ; n7980_not
g34205 not n7971 ; n7971_not
g34206 not n4794 ; n4794_not
g34207 not n9591 ; n9591_not
g34208 not n5766 ; n5766_not
g34209 not n6549 ; n6549_not
g34210 not n5946 ; n5946_not
g34211 not n9636 ; n9636_not
g34212 not n5568 ; n5568_not
g34213 not n9528 ; n9528_not
g34214 not n7584 ; n7584_not
g34215 not n6387 ; n6387_not
g34216 not n9753 ; n9753_not
g34217 not n6765 ; n6765_not
g34218 not n2895 ; n2895_not
g34219 not n2949 ; n2949_not
g34220 not n7593 ; n7593_not
g34221 not n2958 ; n2958_not
g34222 not n7494 ; n7494_not
g34223 not n7386 ; n7386_not
g34224 not n7485 ; n7485_not
g34225 not n4929 ; n4929_not
g34226 not n9690 ; n9690_not
g34227 not n6378 ; n6378_not
g34228 not n3696 ; n3696_not
g34229 not n6747 ; n6747_not
g34230 not n2976 ; n2976_not
g34231 not n2886 ; n2886_not
g34232 not n8286 ; n8286_not
g34233 not n3768 ; n3768_not
g34234 not n8277 ; n8277_not
g34235 not n3759 ; n3759_not
g34236 not n7539 ; n7539_not
g34237 not n8268 ; n8268_not
g34238 not n6783 ; n6783_not
g34239 not n7557 ; n7557_not
g34240 not n7566 ; n7566_not
g34241 not n9519 ; n9519_not
g34242 not n5559 ; n5559_not
g34243 not n8295 ; n8295_not
g34244 not n1779 ; n1779_not
g34245 not n5865 ; n5865_not
g34246 not n5793 ; n5793_not
g34247 not n4668 ; n4668_not
g34248 not n9645 ; n9645_not
g34249 not n7656 ; n7656_not
g34250 not n7647 ; n7647_not
g34251 not n6738 ; n6738_not
g34252 not n6729 ; n6729_not
g34253 not n3795 ; n3795_not
g34254 not n8196 ; n8196_not
g34255 not n3687 ; n3687_not
g34256 not n5667 ; n5667_not
g34257 not n7638 ; n7638_not
g34258 not n6369 ; n6369_not
g34259 not n8187 ; n8187_not
g34260 not n7467 ; n7467_not
g34261 not n5577 ; n5577_not
g34262 not n2868 ; n2868_not
g34263 not n2859 ; n2859_not
g34264 not n8961 ; n8961_not
g34265 not n3678 ; n3678_not
g34266 not n7629 ; n7629_not
g34267 not n7458 ; n7458_not
g34268 not n4677 ; n4677_not
g34269 not n8349 ; n8349_not
g34270 not n9906 ; n9906_not
g34271 not n8970 ; n8970_not
g34272 not n3786 ; n3786_not
g34273 not n2877 ; n2877_not
g34274 not n8178 ; n8178_not
g34275 not n5496 ; n5496_not
g34276 not n4686 ; n4686_not
g34277 not n2994 ; n2994_not
g34278 not n2985 ; n2985_not
g34279 not n9772 ; n9772_not
g34280 not n8926 ; n8926_not
g34281 not n5659 ; n5659_not
g34282 not n8773 ; n8773_not
g34283 not n4858 ; n4858_not
g34284 not n6568 ; n6568_not
g34285 not n9268 ; n9268_not
g34286 not n5884 ; n5884_not
g34287 not n9196 ; n9196_not
g34288 not n6937 ; n6937_not
g34289 not n9187 ; n9187_not
g34290 not n6388 ; n6388_not
g34291 not n6784 ; n6784_not
g34292 not n8737 ; n8737_not
g34293 not n4939 ; n4939_not
g34294 not n9763 ; n9763_not
g34295 not n8962 ; n8962_not
g34296 not n1897 ; n1897_not
g34297 not n9718 ; n9718_not
g34298 not n5668 ; n5668_not
g34299 not n9754 ; n9754_not
g34300 not n9682 ; n9682_not
g34301 not n6298 ; n6298_not
g34302 not n4588 ; n4588_not
g34303 not n8980 ; n8980_not
g34304 not n6487 ; n6487_not
g34305 not n9673 ; n9673_not
g34306 not n6928 ; n6928_not
g34307 not n8971 ; n8971_not
g34308 not n9745 ; n9745_not
g34309 not n8944 ; n8944_not
g34310 not n9259 ; n9259_not
g34311 not n6496 ; n6496_not
g34312 not n4948 ; n4948_not
g34313 not n8755 ; n8755_not
g34314 not n5893 ; n5893_not
g34315 not n4777 ; n4777_not
g34316 not n4795 ; n4795_not
g34317 not n5686 ; n5686_not
g34318 not n6478 ; n6478_not
g34319 not n9826 ; n9826_not
g34320 not n8854 ; n8854_not
g34321 not n1888 ; n1888_not
g34322 not n4786 ; n4786_not
g34323 not n1879 ; n1879_not
g34324 not n8953 ; n8953_not
g34325 not n8935 ; n8935_not
g34326 not n8764 ; n8764_not
g34327 not n4957 ; n4957_not
g34328 not n9628 ; n9628_not
g34329 not n5857 ; n5857_not
g34330 not n6397 ; n6397_not
g34331 not n4894 ; n4894_not
g34332 not n9277 ; n9277_not
g34333 not n8890 ; n8890_not
g34334 not n4966 ; n4966_not
g34335 not n1789 ; n1789_not
g34336 not n6694 ; n6694_not
g34337 not n6739 ; n6739_not
g34338 not n4885 ; n4885_not
g34339 not n6865 ; n6865_not
g34340 not n1996 ; n1996_not
g34341 not n9727 ; n9727_not
g34342 not n9376 ; n9376_not
g34343 not n8674 ; n8674_not
g34344 not n8836 ; n8836_not
g34345 not n9781 ; n9781_not
g34346 not n4678 ; n4678_not
g34347 not n9097 ; n9097_not
g34348 not n9808 ; n9808_not
g34349 not n9691 ; n9691_not
g34350 not n1798 ; n1798_not
g34351 not n4876 ; n4876_not
g34352 not n8827 ; n8827_not
g34353 not n4687 ; n4687_not
g34354 not n8872 ; n8872_not
g34355 not n9295 ; n9295_not
g34356 not n9358 ; n9358_not
g34357 not n8863 ; n8863_not
g34358 not n8548 ; n8548_not
g34359 not n6847 ; n6847_not
g34360 not n4597 ; n4597_not
g34361 not n4984 ; n4984_not
g34362 not n9367 ; n9367_not
g34363 not n9790 ; n9790_not
g34364 not n5875 ; n5875_not
g34365 not n8881 ; n8881_not
g34366 not n8845 ; n8845_not
g34367 not n9088 ; n9088_not
g34368 not n6658 ; n6658_not
g34369 not n9349 ; n9349_not
g34370 not n4759 ; n4759_not
g34371 not n4768 ; n4768_not
g34372 not n8638 ; n8638_not
g34373 not n6586 ; n6586_not
g34374 not n6829 ; n6829_not
g34375 not n5866 ; n5866_not
g34376 not n6775 ; n6775_not
g34377 not n5677 ; n5677_not
g34378 not n8917 ; n8917_not
g34379 not n9385 ; n9385_not
g34380 not n9817 ; n9817_not
g34381 not n9169 ; n9169_not
g34382 not n8782 ; n8782_not
g34383 not n6379 ; n6379_not
g34384 not n9394 ; n9394_not
g34385 not n6577 ; n6577_not
g34386 not n9178 ; n9178_not
g34387 not n1987 ; n1987_not
g34388 not n6883 ; n6883_not
g34389 not n1699 ; n1699_not
g34390 not n6676 ; n6676_not
g34391 not n6667 ; n6667_not
g34392 not n8818 ; n8818_not
g34393 not n1978 ; n1978_not
g34394 not n1969 ; n1969_not
g34395 not n6559 ; n6559_not
g34396 not n6766 ; n6766_not
g34397 not n8908 ; n8908_not
g34398 not n6649 ; n6649_not
g34399 not n6757 ; n6757_not
g34400 not n5578 ; n5578_not
g34401 not n5389 ; n5389_not
g34402 not n5497 ; n5497_not
g34403 not n3985 ; n3985_not
g34404 not n5398 ; n5398_not
g34405 not n3589 ; n3589_not
g34406 not n3598 ; n3598_not
g34407 not n9952 ; n9952_not
g34408 not n9916 ; n9916_not
g34409 not n8494 ; n8494_not
g34410 not n7855 ; n7855_not
g34411 not n2887 ; n2887_not
g34412 not n7819 ; n7819_not
g34413 not n3976 ; n3976_not
g34414 not n9475 ; n9475_not
g34415 not n7792 ; n7792_not
g34416 not n8485 ; n8485_not
g34417 not n9565 ; n9565_not
g34418 not n2878 ; n2878_not
g34419 not n3967 ; n3967_not
g34420 not n7675 ; n7675_not
g34421 not n9943 ; n9943_not
g34422 not n3787 ; n3787_not
g34423 not n7774 ; n7774_not
g34424 not n5767 ; n5767_not
g34425 not n8476 ; n8476_not
g34426 not n9556 ; n9556_not
g34427 not n9484 ; n9484_not
g34428 not n5596 ; n5596_not
g34429 not n9871 ; n9871_not
g34430 not n3499 ; n3499_not
g34431 not n2896 ; n2896_not
g34432 not n8539 ; n8539_not
g34433 not n9574 ; n9574_not
g34434 not n5992 ; n5992_not
g34435 not n7189 ; n7189_not
g34436 not n7198 ; n7198_not
g34437 not n7846 ; n7846_not
g34438 not n8197 ; n8197_not
g34439 not n5587 ; n5587_not
g34440 not n9637 ; n9637_not
g34441 not n5929 ; n5929_not
g34442 not n2698 ; n2698_not
g34443 not n7837 ; n7837_not
g34444 not n9880 ; n9880_not
g34445 not n7909 ; n7909_not
g34446 not n9538 ; n9538_not
g34447 not n3994 ; n3994_not
g34448 not n7828 ; n7828_not
g34449 not n7666 ; n7666_not
g34450 not n7783 ; n7783_not
g34451 not n9466 ; n9466_not
g34452 not n5794 ; n5794_not
g34453 not n8359 ; n8359_not
g34454 not n3868 ; n3868_not
g34455 not n7729 ; n7729_not
g34456 not n5479 ; n5479_not
g34457 not n7369 ; n7369_not
g34458 not n5776 ; n5776_not
g34459 not n7387 ; n7387_not
g34460 not n9493 ; n9493_not
g34461 not n8368 ; n8368_not
g34462 not n8395 ; n8395_not
g34463 not n7693 ; n7693_not
g34464 not n7684 ; n7684_not
g34465 not n2986 ; n2986_not
g34466 not n8386 ; n8386_not
g34467 not n7396 ; n7396_not
g34468 not n9547 ; n9547_not
g34469 not n3697 ; n3697_not
g34470 not n2977 ; n2977_not
g34471 not n3859 ; n3859_not
g34472 not n8377 ; n8377_not
g34473 not n8467 ; n8467_not
g34474 not n3958 ; n3958_not
g34475 not n9925 ; n9925_not
g34476 not n2869 ; n2869_not
g34477 not n3949 ; n3949_not
g34478 not n7468 ; n7468_not
g34479 not n8458 ; n8458_not
g34480 not n7459 ; n7459_not
g34481 not n7279 ; n7279_not
g34482 not n7756 ; n7756_not
g34483 not n8449 ; n8449_not
g34484 not n7099 ; n7099_not
g34485 not n8098 ; n8098_not
g34486 not n7288 ; n7288_not
g34487 not n2797 ; n2797_not
g34488 not n3877 ; n3877_not
g34489 not n9934 ; n9934_not
g34490 not n3886 ; n3886_not
g34491 not n5938 ; n5938_not
g34492 not n7567 ; n7567_not
g34493 not n5488 ; n5488_not
g34494 not n2779 ; n2779_not
g34495 not n5785 ; n5785_not
g34496 not n3895 ; n3895_not
g34497 not n7297 ; n7297_not
g34498 not n8656 ; n8656_not
g34499 not n7954 ; n7954_not
g34500 not n6199 ; n6199_not
g34501 not n3679 ; n3679_not
g34502 not n8647 ; n8647_not
g34503 not n9844 ; n9844_not
g34504 not n5569 ; n5569_not
g34505 not n7963 ; n7963_not
g34506 not n8593 ; n8593_not
g34507 not n9439 ; n9439_not
g34508 not n7576 ; n7576_not
g34509 not n9853 ; n9853_not
g34510 not n9529 ; n9529_not
g34511 not n6991 ; n6991_not
g34512 not n8629 ; n8629_not
g34513 not n7747 ; n7747_not
g34514 not n2599 ; n2599_not
g34515 not n4975 ; n4975_not
g34516 not n2968 ; n2968_not
g34517 not n5983 ; n5983_not
g34518 not n6955 ; n6955_not
g34519 not n7945 ; n7945_not
g34520 not n7927 ; n7927_not
g34521 not n7594 ; n7594_not
g34522 not n9835 ; n9835_not
g34523 not n2959 ; n2959_not
g34524 not n6964 ; n6964_not
g34525 not n6874 ; n6874_not
g34526 not n5965 ; n5965_not
g34527 not n3688 ; n3688_not
g34528 not n7936 ; n7936_not
g34529 not n5974 ; n5974_not
g34530 not n8683 ; n8683_not
g34531 not n5749 ; n5749_not
g34532 not n5695 ; n5695_not
g34533 not n6973 ; n6973_not
g34534 not n8665 ; n8665_not
g34535 not n5758 ; n5758_not
g34536 not n7585 ; n7585_not
g34537 not n7873 ; n7873_not
g34538 not n9862 ; n9862_not
g34539 not n8575 ; n8575_not
g34540 not n3778 ; n3778_not
g34541 not n8179 ; n8179_not
g34542 not n9961 ; n9961_not
g34543 not n7657 ; n7657_not
g34544 not n4579 ; n4579_not
g34545 not n9646 ; n9646_not
g34546 not n4399 ; n4399_not
g34547 not n5299 ; n5299_not
g34548 not n9619 ; n9619_not
g34549 not n7864 ; n7864_not
g34550 not n9286 ; n9286_not
g34551 not n8566 ; n8566_not
g34552 not n8296 ; n8296_not
g34553 not n8557 ; n8557_not
g34554 not n2995 ; n2995_not
g34555 not n9457 ; n9457_not
g34556 not n9655 ; n9655_not
g34557 not n7972 ; n7972_not
g34558 not n9970 ; n9970_not
g34559 not n7558 ; n7558_not
g34560 not n7918 ; n7918_not
g34561 not n9592 ; n9592_not
g34562 not n6838 ; n6838_not
g34563 not n7981 ; n7981_not
g34564 not n7549 ; n7549_not
g34565 not n8269 ; n8269_not
g34566 not n5956 ; n5956_not
g34567 not n4498 ; n4498_not
g34568 not n8188 ; n8188_not
g34569 not n8584 ; n8584_not
g34570 not n8278 ; n8278_not
g34571 not n9664 ; n9664_not
g34572 not n7648 ; n7648_not
g34573 not n8287 ; n8287_not
g34574 not n9448 ; n9448_not
g34575 not n7639 ; n7639_not
g34576 not n7990 ; n7990_not
g34577 not n4489 ; n4489_not
g34578 not n3689 ; n3689_not
g34579 not n7685 ; n7685_not
g34580 not n7658 ; n7658_not
g34581 not n7667 ; n7667_not
g34582 not n2996 ; n2996_not
g34583 not n2978 ; n2978_not
g34584 not n4895 ; n4895_not
g34585 not n5579 ; n5579_not
g34586 not n9737 ; n9737_not
g34587 not n7649 ; n7649_not
g34588 not n9539 ; n9539_not
g34589 not n5588 ; n5588_not
g34590 not n2897 ; n2897_not
g34591 not n4697 ; n4697_not
g34592 not n7676 ; n7676_not
g34593 not n8747 ; n8747_not
g34594 not n8189 ; n8189_not
g34595 not n5786 ; n5786_not
g34596 not n8198 ; n8198_not
g34597 not n2987 ; n2987_not
g34598 not n5876 ; n5876_not
g34599 not n5885 ; n5885_not
g34600 not n7973 ; n7973_not
g34601 not n5984 ; n5984_not
g34602 not n4796 ; n4796_not
g34603 not n7982 ; n7982_not
g34604 not n5957 ; n5957_not
g34605 not n7865 ; n7865_not
g34606 not n9980 ; n9980_not
g34607 not n9269 ; n9269_not
g34608 not n7991 ; n7991_not
g34609 not n9197 ; n9197_not
g34610 not n9971 ; n9971_not
g34611 not n4787 ; n4787_not
g34612 not n9719 ; n9719_not
g34613 not n9188 ; n9188_not
g34614 not n9584 ; n9584_not
g34615 not n9962 ; n9962_not
g34616 not n9953 ; n9953_not
g34617 not n6569 ; n6569_not
g34618 not n7856 ; n7856_not
g34619 not n1898 ; n1898_not
g34620 not n8972 ; n8972_not
g34621 not n5894 ; n5894_not
g34622 not n7892 ; n7892_not
g34623 not n9818 ; n9818_not
g34624 not n4859 ; n4859_not
g34625 not n7919 ; n7919_not
g34626 not n6479 ; n6479_not
g34627 not n5966 ; n5966_not
g34628 not n7928 ; n7928_not
g34629 not n5759 ; n5759_not
g34630 not n9287 ; n9287_not
g34631 not n6488 ; n6488_not
g34632 not n7883 ; n7883_not
g34633 not n8873 ; n8873_not
g34634 not n7946 ; n7946_not
g34635 not n7874 ; n7874_not
g34636 not n6497 ; n6497_not
g34637 not n7955 ; n7955_not
g34638 not n7964 ; n7964_not
g34639 not n9629 ; n9629_not
g34640 not n9593 ; n9593_not
g34641 not n6659 ; n6659_not
g34642 not n9557 ; n9557_not
g34643 not n6668 ; n6668_not
g34644 not n9278 ; n9278_not
g34645 not n9638 ; n9638_not
g34646 not n7766 ; n7766_not
g34647 not n1979 ; n1979_not
g34648 not n7757 ; n7757_not
g34649 not n9935 ; n9935_not
g34650 not n1988 ; n1988_not
g34651 not n6677 ; n6677_not
g34652 not n7595 ; n7595_not
g34653 not n6686 ; n6686_not
g34654 not n7694 ; n7694_not
g34655 not n1997 ; n1997_not
g34656 not n9098 ; n9098_not
g34657 not n9548 ; n9548_not
g34658 not n6695 ; n6695_not
g34659 not n4886 ; n4886_not
g34660 not n9179 ; n9179_not
g34661 not n7748 ; n7748_not
g34662 not n9575 ; n9575_not
g34663 not n7847 ; n7847_not
g34664 not n5993 ; n5993_not
g34665 not n6587 ; n6587_not
g34666 not n7838 ; n7838_not
g34667 not n7829 ; n7829_not
g34668 not n6596 ; n6596_not
g34669 not n4877 ; n4877_not
g34670 not n4778 ; n4778_not
g34671 not n7784 ; n7784_not
g34672 not n9566 ; n9566_not
g34673 not n7793 ; n7793_not
g34674 not n5939 ; n5939_not
g34675 not n3599 ; n3599_not
g34676 not n9944 ; n9944_not
g34677 not n5597 ; n5597_not
g34678 not n7775 ; n7775_not
g34679 not n9674 ; n9674_not
g34680 not n8684 ; n8684_not
g34681 not n9656 ; n9656_not
g34682 not n5399 ; n5399_not
g34683 not n9890 ; n9890_not
g34684 not n8864 ; n8864_not
g34685 not n5678 ; n5678_not
g34686 not n4598 ; n4598_not
g34687 not n5849 ; n5849_not
g34688 not n9881 ; n9881_not
g34689 not n4589 ; n4589_not
g34690 not n3995 ; n3995_not
g34691 not n9467 ; n9467_not
g34692 not n8855 ; n8855_not
g34693 not n9368 ; n9368_not
g34694 not n6857 ; n6857_not
g34695 not n3887 ; n3887_not
g34696 not n4985 ; n4985_not
g34697 not n8765 ; n8765_not
g34698 not n8846 ; n8846_not
g34699 not n2699 ; n2699_not
g34700 not n7199 ; n7199_not
g34701 not n6965 ; n6965_not
g34702 not n8891 ; n8891_not
g34703 not n8477 ; n8477_not
g34704 not n9782 ; n9782_not
g34705 not n4967 ; n4967_not
g34706 not n5858 ; n5858_not
g34707 not n4949 ; n4949_not
g34708 not n9494 ; n9494_not
g34709 not n3968 ; n3968_not
g34710 not n8882 ; n8882_not
g34711 not n9476 ; n9476_not
g34712 not n9791 ; n9791_not
g34713 not n8486 ; n8486_not
g34714 not n3977 ; n3977_not
g34715 not n8495 ; n8495_not
g34716 not n6848 ; n6848_not
g34717 not n8756 ; n8756_not
g34718 not n9359 ; n9359_not
g34719 not n6893 ; n6893_not
g34720 not n8585 ; n8585_not
g34721 not n6974 ; n6974_not
g34722 not n8648 ; n8648_not
g34723 not n9377 ; n9377_not
g34724 not n4994 ; n4994_not
g34725 not n8774 ; n8774_not
g34726 not n9449 ; n9449_not
g34727 not n9395 ; n9395_not
g34728 not n8639 ; n8639_not
g34729 not n4499 ; n4499_not
g34730 not n6749 ; n6749_not
g34731 not n9386 ; n9386_not
g34732 not n9845 ; n9845_not
g34733 not n9854 ; n9854_not
g34734 not n9692 ; n9692_not
g34735 not n8792 ; n8792_not
g34736 not n8783 ; n8783_not
g34737 not n6299 ; n6299_not
g34738 not n9872 ; n9872_not
g34739 not n6866 ; n6866_not
g34740 not n9458 ; n9458_not
g34741 not n8837 ; n8837_not
g34742 not n6938 ; n6938_not
g34743 not n8657 ; n8657_not
g34744 not n8549 ; n8549_not
g34745 not n6956 ; n6956_not
g34746 not n9863 ; n9863_not
g34747 not n8558 ; n8558_not
g34748 not n8567 ; n8567_not
g34749 not n9809 ; n9809_not
g34750 not n8675 ; n8675_not
g34751 not n6884 ; n6884_not
g34752 not n8576 ; n8576_not
g34753 not n6776 ; n6776_not
g34754 not n8297 ; n8297_not
g34755 not n6947 ; n6947_not
g34756 not n8990 ; n8990_not
g34757 not n8738 ; n8738_not
g34758 not n8936 ; n8936_not
g34759 not n9755 ; n9755_not
g34760 not n8981 ; n8981_not
g34761 not n7487 ; n7487_not
g34762 not n2879 ; n2879_not
g34763 not n4976 ; n4976_not
g34764 not n2888 ; n2888_not
g34765 not n5498 ; n5498_not
g34766 not n8378 ; n8378_not
g34767 not n7478 ; n7478_not
g34768 not n9827 ; n9827_not
g34769 not n8945 ; n8945_not
g34770 not n7469 ; n7469_not
g34771 not n2798 ; n2798_not
g34772 not n3698 ; n3698_not
g34773 not n6758 ; n6758_not
g34774 not n6767 ; n6767_not
g34775 not n6398 ; n6398_not
g34776 not n8729 ; n8729_not
g34777 not n7388 ; n7388_not
g34778 not n7577 ; n7577_not
g34779 not n7568 ; n7568_not
g34780 not n8279 ; n8279_not
g34781 not n6389 ; n6389_not
g34782 not n8288 ; n8288_not
g34783 not n3779 ; n3779_not
g34784 not n6785 ; n6785_not
g34785 not n5768 ; n5768_not
g34786 not n9665 ; n9665_not
g34787 not n9746 ; n9746_not
g34788 not n8387 ; n8387_not
g34789 not n8918 ; n8918_not
g34790 not n8927 ; n8927_not
g34791 not n9836 ; n9836_not
g34792 not n3869 ; n3869_not
g34793 not n9773 ; n9773_not
g34794 not n3878 ; n3878_not
g34795 not n2789 ; n2789_not
g34796 not n3896 ; n3896_not
g34797 not n9485 ; n9485_not
g34798 not n7289 ; n7289_not
g34799 not n8909 ; n8909_not
g34800 not n6839 ; n6839_not
g34801 not n8459 ; n8459_not
g34802 not n9764 ; n9764_not
g34803 not n9728 ; n9728_not
g34804 not n3959 ; n3959_not
g34805 not n8468 ; n8468_not
g34806 not n3797 ; n3797_not
g34807 not n9683 ; n9683_not
g34808 not n8369 ; n8369_not
g34809 not n8954 ; n8954_not
g34810 not n6794 ; n6794_not
g34811 not n5687 ; n5687_not
g34812 not n6929 ; n6929_not
g34813 not n7397 ; n7397_not
g34814 not n4958 ; n4958_not
g34815 not n8396 ; n8396_not
g34816 not n6875 ; n6875_not
g34817 not n9657 ; n9657_not
g34818 not n5985 ; n5985_not
g34819 not n9477 ; n9477_not
g34820 not n9396 ; n9396_not
g34821 not n5958 ; n5958_not
g34822 not n9567 ; n9567_not
g34823 not n9558 ; n9558_not
g34824 not n4878 ; n4878_not
g34825 not n8982 ; n8982_not
g34826 not n9279 ; n9279_not
g34827 not n4959 ; n4959_not
g34828 not n5589 ; n5589_not
g34829 not n8964 ; n8964_not
g34830 not n9549 ; n9549_not
g34831 not n9495 ; n9495_not
g34832 not n9189 ; n9189_not
g34833 not n9459 ; n9459_not
g34834 not n9684 ; n9684_not
g34835 not n5499 ; n5499_not
g34836 not a[0] ; a[0]_not
g34837 not n5787 ; n5787_not
g34838 not n9198 ; n9198_not
g34839 not n5796 ; n5796_not
g34840 not n4896 ; n4896_not
g34841 not n4887 ; n4887_not
g34842 not n6399 ; n6399_not
g34843 not n9675 ; n9675_not
g34844 not n9594 ; n9594_not
g34845 not n4995 ; n4995_not
g34846 not n9387 ; n9387_not
g34847 not n5994 ; n5994_not
g34848 not n5949 ; n5949_not
g34849 not n9378 ; n9378_not
g34850 not n9585 ; n9585_not
g34851 not n4869 ; n4869_not
g34852 not n9288 ; n9288_not
g34853 not n4986 ; n4986_not
g34854 not n9468 ; n9468_not
g34855 not n4977 ; n4977_not
g34856 not n9639 ; n9639_not
g34857 not n8676 ; n8676_not
g34858 not n7668 ; n7668_not
g34859 not n8775 ; n8775_not
g34860 not n7659 ; n7659_not
g34861 not n8766 ; n8766_not
g34862 not n8757 ; n8757_not
g34863 not n8748 ; n8748_not
g34864 not n8739 ; n8739_not
g34865 not n5688 ; n5688_not
g34866 not n2988 ; n2988_not
g34867 not n8199 ; n8199_not
g34868 not n6939 ; n6939_not
g34869 not n6948 ; n6948_not
g34870 not n9918 ; n9918_not
g34871 not n9972 ; n9972_not
g34872 not n2979 ; n2979_not
g34873 not n6957 ; n6957_not
g34874 not n9576 ; n9576_not
g34875 not n7596 ; n7596_not
g34876 not n9837 ; n9837_not
g34877 not n8694 ; n8694_not
g34878 not n7578 ; n7578_not
g34879 not n8685 ; n8685_not
g34880 not n9828 ; n9828_not
g34881 not n6966 ; n6966_not
g34882 not n8469 ; n8469_not
g34883 not n7767 ; n7767_not
g34884 not n8874 ; n8874_not
g34885 not n9792 ; n9792_not
g34886 not n9693 ; n9693_not
g34887 not n7758 ; n7758_not
g34888 not n8856 ; n8856_not
g34889 not n8649 ; n8649_not
g34890 not n6858 ; n6858_not
g34891 not n7749 ; n7749_not
g34892 not n8847 ; n8847_not
g34893 not n5778 ; n5778_not
g34894 not n8838 ; n8838_not
g34895 not n6876 ; n6876_not
g34896 not n6885 ; n6885_not
g34897 not n7686 ; n7686_not
g34898 not n6894 ; n6894_not
g34899 not n5679 ; n5679_not
g34900 not n8793 ; n8793_not
g34901 not n9819 ; n9819_not
g34902 not n2997 ; n2997_not
g34903 not n8784 ; n8784_not
g34904 not n9864 ; n9864_not
g34905 not n9909 ; n9909_not
g34906 not n7677 ; n7677_not
g34907 not n9873 ; n9873_not
g34908 not n3798 ; n3798_not
g34909 not n9882 ; n9882_not
g34910 not n8379 ; n8379_not
g34911 not n8496 ; n8496_not
g34912 not n3978 ; n3978_not
g34913 not n7398 ; n7398_not
g34914 not n8487 ; n8487_not
g34915 not n9891 ; n9891_not
g34916 not n3969 ; n3969_not
g34917 not n7389 ; n7389_not
g34918 not n8478 ; n8478_not
g34919 not n8397 ; n8397_not
g34920 not n3897 ; n3897_not
g34921 not n8388 ; n8388_not
g34922 not n3888 ; n3888_not
g34923 not n2799 ; n2799_not
g34924 not n7569 ; n7569_not
g34925 not n6678 ; n6678_not
g34926 not n8289 ; n8289_not
g34927 not n8658 ; n8658_not
g34928 not n6975 ; n6975_not
g34929 not n6984 ; n6984_not
g34930 not n8586 ; n8586_not
g34931 not n9846 ; n9846_not
g34932 not n2898 ; n2898_not
g34933 not n8298 ; n8298_not
g34934 not n6993 ; n6993_not
g34935 not n9666 ; n9666_not
g34936 not n6849 ; n6849_not
g34937 not n8595 ; n8595_not
g34938 not n9855 ; n9855_not
g34939 not n7497 ; n7497_not
g34940 not n7488 ; n7488_not
g34941 not n2889 ; n2889_not
g34942 not n7479 ; n7479_not
g34943 not n8577 ; n8577_not
g34944 not n8568 ; n8568_not
g34945 not n4698 ; n4698_not
g34946 not n7965 ; n7965_not
g34947 not n1899 ; n1899_not
g34948 not n9738 ; n9738_not
g34949 not n7974 ; n7974_not
g34950 not n7983 ; n7983_not
g34951 not n7866 ; n7866_not
g34952 not n6759 ; n6759_not
g34953 not n5868 ; n5868_not
g34954 not n6768 ; n6768_not
g34955 not n9981 ; n9981_not
g34956 not n7992 ; n7992_not
g34957 not n6777 ; n6777_not
g34958 not n6786 ; n6786_not
g34959 not n9747 ; n9747_not
g34960 not n9963 ; n9963_not
g34961 not n8991 ; n8991_not
g34962 not n5895 ; n5895_not
g34963 not n8892 ; n8892_not
g34964 not n6498 ; n6498_not
g34965 not n9783 ; n9783_not
g34966 not n7893 ; n7893_not
g34967 not n4797 ; n4797_not
g34968 not n7929 ; n7929_not
g34969 not n4788 ; n4788_not
g34970 not n6588 ; n6588_not
g34971 not n7884 ; n7884_not
g34972 not n7875 ; n7875_not
g34973 not n6669 ; n6669_not
g34974 not n1989 ; n1989_not
g34975 not n7947 ; n7947_not
g34976 not n6687 ; n6687_not
g34977 not n9099 ; n9099_not
g34978 not n6696 ; n6696_not
g34979 not n5877 ; n5877_not
g34980 not n7848 ; n7848_not
g34981 not n5859 ; n5859_not
g34982 not n7839 ; n7839_not
g34983 not n8955 ; n8955_not
g34984 not n5769 ; n5769_not
g34985 not n8946 ; n8946_not
g34986 not n9765 ; n9765_not
g34987 not n6795 ; n6795_not
g34988 not n9954 ; n9954_not
g34989 not n7794 ; n7794_not
g34990 not n8928 ; n8928_not
g34991 not n8919 ; n8919_not
g34992 not n9774 ; n9774_not
g34993 not n4599 ; n4599_not
g34994 not n7785 ; n7785_not
g34995 not n9936 ; n9936_not
g34996 not n8883 ; n8883_not
g34997 not n9756 ; n9756_not
g34998 not n9729 ; n9729_not
g34999 not n7857 ; n7857_not
g35000 not n8973 ; n8973_not
g35001 not n7885 ; n7885_not
g35002 not n5797 ; n5797_not
g35003 not n9586 ; n9586_not
g35004 not n9649 ; n9649_not
g35005 not n7939 ; n7939_not
g35006 not n3799 ; n3799_not
g35007 not n7876 ; n7876_not
g35008 not n7993 ; n7993_not
g35009 not n5977 ; n5977_not
g35010 not n7579 ; n7579_not
g35011 not n7597 ; n7597_not
g35012 not n7795 ; n7795_not
g35013 not n7588 ; n7588_not
g35014 not b[0] ; b[0]_not
g35015 not n9577 ; n9577_not
g35016 not n9496 ; n9496_not
g35017 not n2989 ; n2989_not
g35018 not n5599 ; n5599_not
g35019 not n9973 ; n9973_not
g35020 not n8389 ; n8389_not
g35021 not n9883 ; n9883_not
g35022 not n8398 ; n8398_not
g35023 not n9937 ; n9937_not
g35024 not n7768 ; n7768_not
g35025 not n8974 ; n8974_not
g35026 not n9919 ; n9919_not
g35027 not n2998 ; n2998_not
g35028 not n5788 ; n5788_not
g35029 not n9559 ; n9559_not
g35030 not n7759 ; n7759_not
g35031 not n7399 ; n7399_not
g35032 not n7498 ; n7498_not
g35033 not n2899 ; n2899_not
g35034 not n9595 ; n9595_not
g35035 not n9982 ; n9982_not
g35036 not n7867 ; n7867_not
g35037 not n7489 ; n7489_not
g35038 not n7984 ; n7984_not
g35039 not n7849 ; n7849_not
g35040 not n7894 ; n7894_not
g35041 not n7687 ; n7687_not
g35042 not n5959 ; n5959_not
g35043 not n9568 ; n9568_not
g35044 not n7948 ; n7948_not
g35045 not n7858 ; n7858_not
g35046 not n9847 ; n9847_not
g35047 not n9928 ; n9928_not
g35048 not n7678 ; n7678_not
g35049 not n5986 ; n5986_not
g35050 not n8299 ; n8299_not
g35051 not n9748 ; n9748_not
g35052 not n6787 ; n6787_not
g35053 not n8992 ; n8992_not
g35054 not n9757 ; n9757_not
g35055 not a[1] ; a[1]_not
g35056 not n8947 ; n8947_not
g35057 not n8965 ; n8965_not
g35058 not n8956 ; n8956_not
g35059 not n9766 ; n9766_not
g35060 not n6796 ; n6796_not
g35061 not n8938 ; n8938_not
g35062 not n6877 ; n6877_not
g35063 not n9676 ; n9676_not
g35064 not n8839 ; n8839_not
g35065 not n6859 ; n6859_not
g35066 not n4798 ; n4798_not
g35067 not n8848 ; n8848_not
g35068 not n6697 ; n6697_not
g35069 not n8857 ; n8857_not
g35070 not n9793 ; n9793_not
g35071 not n4978 ; n4978_not
g35072 not n8875 ; n8875_not
g35073 not n9784 ; n9784_not
g35074 not n8893 ; n8893_not
g35075 not n9775 ; n9775_not
g35076 not n8929 ; n8929_not
g35077 not n9397 ; n9397_not
g35078 not n6499 ; n6499_not
g35079 not n5887 ; n5887_not
g35080 not n9199 ; n9199_not
g35081 not n4789 ; n4789_not
g35082 not n6589 ; n6589_not
g35083 not n5878 ; n5878_not
g35084 not n4879 ; n4879_not
g35085 not n8983 ; n8983_not
g35086 not n6679 ; n6679_not
g35087 not n6688 ; n6688_not
g35088 not n5896 ; n5896_not
g35089 not n4888 ; n4888_not
g35090 not n6778 ; n6778_not
g35091 not n6769 ; n6769_not
g35092 not n5869 ; n5869_not
g35093 not n8776 ; n8776_not
g35094 not n8767 ; n8767_not
g35095 not n1999 ; n1999_not
g35096 not n4897 ; n4897_not
g35097 not n9694 ; n9694_not
g35098 not n9739 ; n9739_not
g35099 not n9298 ; n9298_not
g35100 not n9289 ; n9289_not
g35101 not n4699 ; n4699_not
g35102 not n8677 ; n8677_not
g35103 not n6967 ; n6967_not
g35104 not n8668 ; n8668_not
g35105 not n9658 ; n9658_not
g35106 not n8659 ; n8659_not
g35107 not n6976 ; n6976_not
g35108 not n6985 ; n6985_not
g35109 not n9667 ; n9667_not
g35110 not n6994 ; n6994_not
g35111 not n5698 ; n5698_not
g35112 not n5995 ; n5995_not
g35113 not n8596 ; n8596_not
g35114 not n9856 ; n9856_not
g35115 not n8587 ; n8587_not
g35116 not n9892 ; n9892_not
g35117 not n3889 ; n3889_not
g35118 not n9478 ; n9478_not
g35119 not n8479 ; n8479_not
g35120 not n8488 ; n8488_not
g35121 not n3979 ; n3979_not
g35122 not n3988 ; n3988_not
g35123 not n8497 ; n8497_not
g35124 not n3997 ; n3997_not
g35125 not n9874 ; n9874_not
g35126 not n6598 ; n6598_not
g35127 not n8569 ; n8569_not
g35128 not n8749 ; n8749_not
g35129 not n8785 ; n8785_not
g35130 not n5689 ; n5689_not
g35131 not n4996 ; n4996_not
g35132 not n8794 ; n8794_not
g35133 not n9829 ; n9829_not
g35134 not n4987 ; n4987_not
g35135 not n6895 ; n6895_not
g35136 not n6949 ; n6949_not
g35137 not n5968 ; n5968_not
g35138 not n8686 ; n8686_not
g35139 not n9838 ; n9838_not
g35140 not n8695 ; n8695_not
g35141 not n6886 ; n6886_not
g35142 not n6958 ; n6958_not
g35143 not n5879 ; n5879_not
g35144 not b[1] ; b[1]_not
g35145 not n5888 ; n5888_not
g35146 not n9785 ; n9785_not
g35147 not n9929 ; n9929_not
g35148 not n5798 ; n5798_not
g35149 not n9893 ; n9893_not
g35150 not a[2] ; a[2]_not
g35151 not n9677 ; n9677_not
g35152 not n5699 ; n5699_not
g35153 not n9758 ; n9758_not
g35154 not n9839 ; n9839_not
g35155 not n9956 ; n9956_not
g35156 not n9767 ; n9767_not
g35157 not n9974 ; n9974_not
g35158 not n9848 ; n9848_not
g35159 not n9776 ; n9776_not
g35160 not n9947 ; n9947_not
g35161 not n5897 ; n5897_not
g35162 not n9695 ; n9695_not
g35163 not n9983 ; n9983_not
g35164 not n9938 ; n9938_not
g35165 not n9992 ; n9992_not
g35166 not n5789 ; n5789_not
g35167 not n9866 ; n9866_not
g35168 not n9668 ; n9668_not
g35169 not n9875 ; n9875_not
g35170 not n6977 ; n6977_not
g35171 not n8498 ; n8498_not
g35172 not n3989 ; n3989_not
g35173 not n3998 ; n3998_not
g35174 not n6968 ; n6968_not
g35175 not n4799 ; n4799_not
g35176 not n8588 ; n8588_not
g35177 not n6599 ; n6599_not
g35178 not n8597 ; n8597_not
g35179 not n6698 ; n6698_not
g35180 not n6986 ; n6986_not
g35181 not n8669 ; n8669_not
g35182 not n7769 ; n7769_not
g35183 not n7697 ; n7697_not
g35184 not n7688 ; n7688_not
g35185 not n7679 ; n7679_not
g35186 not n2999 ; n2999_not
g35187 not n7598 ; n7598_not
g35188 not n7589 ; n7589_not
g35189 not n7499 ; n7499_not
g35190 not n4898 ; n4898_not
g35191 not n8399 ; n8399_not
g35192 not n9299 ; n9299_not
g35193 not n4889 ; n4889_not
g35194 not n6995 ; n6995_not
g35195 not n8975 ; n8975_not
g35196 not n8786 ; n8786_not
g35197 not n8966 ; n8966_not
g35198 not n6896 ; n6896_not
g35199 not n8957 ; n8957_not
g35200 not n8948 ; n8948_not
g35201 not n6878 ; n6878_not
g35202 not n8939 ; n8939_not
g35203 not n6797 ; n6797_not
g35204 not n6869 ; n6869_not
g35205 not n8849 ; n8849_not
g35206 not n8858 ; n8858_not
g35207 not n8867 ; n8867_not
g35208 not n8876 ; n8876_not
g35209 not n8894 ; n8894_not
g35210 not n8678 ; n8678_not
g35211 not n8696 ; n8696_not
g35212 not n6959 ; n6959_not
g35213 not n6887 ; n6887_not
g35214 not n6779 ; n6779_not
g35215 not n8768 ; n8768_not
g35216 not n8993 ; n8993_not
g35217 not n8984 ; n8984_not
g35218 not n8777 ; n8777_not
g35219 not n8687 ; n8687_not
g35220 not n6788 ; n6788_not
g35221 not n8795 ; n8795_not
g35222 not n7985 ; n7985_not
g35223 not n7895 ; n7895_not
g35224 not n4988 ; n4988_not
g35225 not n7994 ; n7994_not
g35226 not n7877 ; n7877_not
g35227 not n9596 ; n9596_not
g35228 not n9488 ; n9488_not
g35229 not n5996 ; n5996_not
g35230 not n9578 ; n9578_not
g35231 not n9569 ; n9569_not
g35232 not n7886 ; n7886_not
g35233 not n9479 ; n9479_not
g35234 not n7949 ; n7949_not
g35235 not n7958 ; n7958_not
g35236 not n9587 ; n9587_not
g35237 not n7868 ; n7868_not
g35238 not n7967 ; n7967_not
g35239 not n4979 ; n4979_not
g35240 not n7778 ; n7778_not
g35241 not n4997 ; n4997_not
g35242 not n5969 ; n5969_not
g35243 not n9398 ; n9398_not
g35244 not n7796 ; n7796_not
g35245 not n9497 ; n9497_not
g35246 not n5978 ; n5978_not
g35247 not n7859 ; n7859_not
g35248 not n7959 ; n7959_not
g35249 not n8949 ; n8949_not
g35250 not n7869 ; n7869_not
g35251 not n8769 ; n8769_not
g35252 not n9849 ; n9849_not
g35253 not n8688 ; n8688_not
g35254 not n7896 ; n7896_not
g35255 not n9786 ; n9786_not
g35256 not n8886 ; n8886_not
g35257 not n8877 ; n8877_not
g35258 not b[2] ; b[2]_not
g35259 not n8868 ; n8868_not
g35260 not n9795 ; n9795_not
g35261 not n8859 ; n8859_not
g35262 not n9777 ; n9777_not
g35263 not n7887 ; n7887_not
g35264 not n6888 ; n6888_not
g35265 not n6897 ; n6897_not
g35266 not n7878 ; n7878_not
g35267 not n8796 ; n8796_not
g35268 not n8787 ; n8787_not
g35269 not n3999 ; n3999_not
g35270 not n9876 ; n9876_not
g35271 not n7995 ; n7995_not
g35272 not n9885 ; n9885_not
g35273 not n8499 ; n8499_not
g35274 not n9966 ; n9966_not
g35275 not n9957 ; n9957_not
g35276 not n9894 ; n9894_not
g35277 not n7986 ; n7986_not
g35278 not n7797 ; n7797_not
g35279 not n9948 ; n9948_not
g35280 not n7788 ; n7788_not
g35281 not n7779 ; n7779_not
g35282 not n9939 ; n9939_not
g35283 not n7689 ; n7689_not
g35284 not n7698 ; n7698_not
g35285 not n9597 ; n9597_not
g35286 not n9858 ; n9858_not
g35287 not n8697 ; n8697_not
g35288 not n7968 ; n7968_not
g35289 not n8679 ; n8679_not
g35290 not n7977 ; n7977_not
g35291 not n6969 ; n6969_not
g35292 not n9993 ; n9993_not
g35293 not n9678 ; n9678_not
g35294 not n9975 ; n9975_not
g35295 not n6987 ; n6987_not
g35296 not n6978 ; n6978_not
g35297 not n6996 ; n6996_not
g35298 not n8589 ; n8589_not
g35299 not n5799 ; n5799_not
g35300 not a[3] ; a[3]_not
g35301 not n9867 ; n9867_not
g35302 not n9498 ; n9498_not
g35303 not n9588 ; n9588_not
g35304 not n5979 ; n5979_not
g35305 not n6789 ; n6789_not
g35306 not n9669 ; n9669_not
g35307 not n8994 ; n8994_not
g35308 not n6699 ; n6699_not
g35309 not n9489 ; n9489_not
g35310 not n6798 ; n6798_not
g35311 not n9399 ; n9399_not
g35312 not n8958 ; n8958_not
g35313 not n8985 ; n8985_not
g35314 not n5889 ; n5889_not
g35315 not n8967 ; n8967_not
g35316 not n5898 ; n5898_not
g35317 not n8895 ; n8895_not
g35318 not n9687 ; n9687_not
g35319 not n4899 ; n4899_not
g35320 not n5997 ; n5997_not
g35321 not n4989 ; n4989_not
g35322 not n9579 ; n9579_not
g35323 not n4998 ; n4998_not
g35324 not n9696 ; n9696_not
g35325 not n7969 ; n7969_not
g35326 not n9994 ; n9994_not
g35327 not n8689 ; n8689_not
g35328 not n7978 ; n7978_not
g35329 not n9859 ; n9859_not
g35330 not n6997 ; n6997_not
g35331 not n9985 ; n9985_not
g35332 not n6988 ; n6988_not
g35333 not b[3] ; b[3]_not
g35334 not n9499 ; n9499_not
g35335 not n6979 ; n6979_not
g35336 not n9688 ; n9688_not
g35337 not n7699 ; n7699_not
g35338 not n5899 ; n5899_not
g35339 not n9679 ; n9679_not
g35340 not n7789 ; n7789_not
g35341 not n9949 ; n9949_not
g35342 not n7798 ; n7798_not
g35343 not n9895 ; n9895_not
g35344 not n9886 ; n9886_not
g35345 not n9967 ; n9967_not
g35346 not n4999 ; n4999_not
g35347 not n9877 ; n9877_not
g35348 not n9976 ; n9976_not
g35349 not n9868 ; n9868_not
g35350 not a[4] ; a[4]_not
g35351 not n8995 ; n8995_not
g35352 not n7987 ; n7987_not
g35353 not n8779 ; n8779_not
g35354 not n8788 ; n8788_not
g35355 not n9589 ; n9589_not
g35356 not n8977 ; n8977_not
g35357 not n8797 ; n8797_not
g35358 not n5989 ; n5989_not
g35359 not n8959 ; n8959_not
g35360 not n6889 ; n6889_not
g35361 not n7888 ; n7888_not
g35362 not n6799 ; n6799_not
g35363 not n9796 ; n9796_not
g35364 not n8869 ; n8869_not
g35365 not n9778 ; n9778_not
g35366 not n8878 ; n8878_not
g35367 not n7897 ; n7897_not
g35368 not n8896 ; n8896_not
g35369 not n8887 ; n8887_not
g35370 not n6898 ; n6898_not
g35371 not n5998 ; n5998_not
g35372 not n8986 ; n8986_not
g35373 not n9958 ; n9958_not
g35374 not n8698 ; n8698_not
g35375 not n7879 ; n7879_not
g35376 not n8897 ; n8897_not
g35377 not n9896 ; n9896_not
g35378 not n9797 ; n9797_not
g35379 not n9779 ; n9779_not
g35380 not n7799 ; n7799_not
g35381 not n7898 ; n7898_not
g35382 not n9959 ; n9959_not
g35383 not n9599 ; n9599_not
g35384 not n7889 ; n7889_not
g35385 not n9995 ; n9995_not
g35386 not b[4] ; b[4]_not
g35387 not n8996 ; n8996_not
g35388 not a[5] ; a[5]_not
g35389 not n9788 ; n9788_not
g35390 not n8879 ; n8879_not
g35391 not n9986 ; n9986_not
g35392 not n7997 ; n7997_not
g35393 not n8888 ; n8888_not
g35394 not n9689 ; n9689_not
g35395 not n6998 ; n6998_not
g35396 not n8798 ; n8798_not
g35397 not n7979 ; n7979_not
g35398 not n8789 ; n8789_not
g35399 not n8978 ; n8978_not
g35400 not n9968 ; n9968_not
g35401 not n6989 ; n6989_not
g35402 not n9977 ; n9977_not
g35403 not n9887 ; n9887_not
g35404 not n6899 ; n6899_not
g35405 not n9878 ; n9878_not
g35406 not n8699 ; n8699_not
g35407 not n7989 ; n7989_not
g35408 not n9969 ; n9969_not
g35409 not a[6] ; a[6]_not
g35410 not b[5] ; b[5]_not
g35411 not n9978 ; n9978_not
g35412 not n9987 ; n9987_not
g35413 not n9996 ; n9996_not
g35414 not n7899 ; n7899_not
g35415 not n7998 ; n7998_not
g35416 not n9798 ; n9798_not
g35417 not n9879 ; n9879_not
g35418 not n8997 ; n8997_not
g35419 not n6999 ; n6999_not
g35420 not n8898 ; n8898_not
g35421 not n9897 ; n9897_not
g35422 not n8799 ; n8799_not
g35423 not n9699 ; n9699_not
g35424 not n8979 ; n8979_not
g35425 not n9789 ; n9789_not
g35426 not n8889 ; n8889_not
g35427 not n9898 ; n9898_not
g35428 not n7999 ; n7999_not
g35429 not a[7] ; a[7]_not
g35430 not n8989 ; n8989_not
g35431 not n8998 ; n8998_not
g35432 not n9799 ; n9799_not
g35433 not b[6] ; b[6]_not
g35434 not n9997 ; n9997_not
g35435 not n8899 ; n8899_not
g35436 not n9988 ; n9988_not
g35437 not n9979 ; n9979_not
g35438 not a[8] ; a[8]_not
g35439 not b[7] ; b[7]_not
g35440 not n9989 ; n9989_not
g35441 not n9899 ; n9899_not
g35442 not n8999 ; n8999_not
g35443 not n9998 ; n9998_not
g35444 not b[8] ; b[8]_not
g35445 not a[9] ; a[9]_not
g35446 not n9999 ; n9999_not
g35447 not b[9] ; b[9]_not
g35448 not n10000 ; n10000_not
g35449 not n10010 ; n10010_not
g35450 not n10001 ; n10001_not
g35451 not n11000 ; n11000_not
g35452 not n10100 ; n10100_not
g35453 not n20000 ; n20000_not
g35454 not n10011 ; n10011_not
g35455 not n10110 ; n10110_not
g35456 not n20010 ; n20010_not
g35457 not n11001 ; n11001_not
g35458 not n20100 ; n20100_not
g35459 not n12000 ; n12000_not
g35460 not n21000 ; n21000_not
g35461 not n10002 ; n10002_not
g35462 not n20001 ; n20001_not
g35463 not n10101 ; n10101_not
g35464 not n10020 ; n10020_not
g35465 not n11010 ; n11010_not
g35466 not n10200 ; n10200_not
g35467 not n10003 ; n10003_not
g35468 not n20020 ; n20020_not
g35469 not n20101 ; n20101_not
g35470 not n10111 ; n10111_not
g35471 not n10012 ; n10012_not
g35472 not n20011 ; n20011_not
g35473 not n10120 ; n10120_not
g35474 not n20110 ; n20110_not
g35475 not n10102 ; n10102_not
g35476 not n10021 ; n10021_not
g35477 not n10030 ; n10030_not
g35478 not n10300 ; n10300_not
g35479 not n10201 ; n10201_not
g35480 not n10210 ; n10210_not
g35481 not n21001 ; n21001_not
g35482 not n21010 ; n21010_not
g35483 not n20200 ; n20200_not
g35484 not n11020 ; n11020_not
g35485 not n13000 ; n13000_not
g35486 not n12010 ; n12010_not
g35487 not n11002 ; n11002_not
g35488 not n11101 ; n11101_not
g35489 not n21100 ; n21100_not
g35490 not n12100 ; n12100_not
g35491 not n11200 ; n11200_not
g35492 not n22000 ; n22000_not
g35493 not n11011 ; n11011_not
g35494 not n20002 ; n20002_not
g35495 not n11110 ; n11110_not
g35496 not n21011 ; n21011_not
g35497 not n21020 ; n21020_not
g35498 not n23000 ; n23000_not
g35499 not n10031 ; n10031_not
g35500 not n12020 ; n12020_not
g35501 not n10202 ; n10202_not
g35502 not n20102 ; n20102_not
g35503 not n12200 ; n12200_not
g35504 not n13100 ; n13100_not
g35505 not n12110 ; n12110_not
g35506 not n21101 ; n21101_not
g35507 not n21110 ; n21110_not
g35508 not n13010 ; n13010_not
g35509 not n13001 ; n13001_not
g35510 not n10112 ; n10112_not
g35511 not n10121 ; n10121_not
g35512 not n12101 ; n12101_not
g35513 not n10130 ; n10130_not
g35514 not n10103 ; n10103_not
g35515 not n11030 ; n11030_not
g35516 not n20120 ; n20120_not
g35517 not n14000 ; n14000_not
g35518 not n11102 ; n11102_not
g35519 not n11111 ; n11111_not
g35520 not n11120 ; n11120_not
g35521 not n22001 ; n22001_not
g35522 not n20012 ; n20012_not
g35523 not n11201 ; n11201_not
g35524 not n20021 ; n20021_not
g35525 not n11210 ; n11210_not
g35526 not n10400 ; n10400_not
g35527 not n12011 ; n12011_not
g35528 not n10220 ; n10220_not
g35529 not n20210 ; n20210_not
g35530 not n12002 ; n12002_not
g35531 not n20201 ; n20201_not
g35532 not n20003 ; n20003_not
g35533 not n20030 ; n20030_not
g35534 not n11021 ; n11021_not
g35535 not n22100 ; n22100_not
g35536 not n22010 ; n22010_not
g35537 not n10301 ; n10301_not
g35538 not n20300 ; n20300_not
g35539 not n10004 ; n10004_not
g35540 not n21002 ; n21002_not
g35541 not n10040 ; n10040_not
g35542 not n10022 ; n10022_not
g35543 not n10013 ; n10013_not
g35544 not n11202 ; n11202_not
g35545 not n23001 ; n23001_not
g35546 not n11211 ; n11211_not
g35547 not n12003 ; n12003_not
g35548 not n11220 ; n11220_not
g35549 not n10050 ; n10050_not
g35550 not n10320 ; n10320_not
g35551 not n21030 ; n21030_not
g35552 not n22110 ; n22110_not
g35553 not n13110 ; n13110_not
g35554 not n22002 ; n22002_not
g35555 not n20400 ; n20400_not
g35556 not n11121 ; n11121_not
g35557 not n11301 ; n11301_not
g35558 not n13101 ; n13101_not
g35559 not n12012 ; n12012_not
g35560 not n21300 ; n21300_not
g35561 not n12300 ; n12300_not
g35562 not n10014 ; n10014_not
g35563 not n10005 ; n10005_not
g35564 not n21003 ; n21003_not
g35565 not n20013 ; n20013_not
g35566 not n12021 ; n12021_not
g35567 not n12030 ; n12030_not
g35568 not n20310 ; n20310_not
g35569 not n21201 ; n21201_not
g35570 not n20220 ; n20220_not
g35571 not n20112 ; n20112_not
g35572 not n14100 ; n14100_not
g35573 not n20121 ; n20121_not
g35574 not n11400 ; n11400_not
g35575 not n10041 ; n10041_not
g35576 not n10221 ; n10221_not
g35577 not n13020 ; n13020_not
g35578 not n20130 ; n20130_not
g35579 not n21111 ; n21111_not
g35580 not n13011 ; n13011_not
g35581 not n14010 ; n14010_not
g35582 not n21120 ; n21120_not
g35583 not n14001 ; n14001_not
g35584 not n10311 ; n10311_not
g35585 not n22020 ; n22020_not
g35586 not n11310 ; n11310_not
g35587 not n10302 ; n10302_not
g35588 not n20103 ; n20103_not
g35589 not n20004 ; n20004_not
g35590 not n23100 ; n23100_not
g35591 not n10032 ; n10032_not
g35592 not n10203 ; n10203_not
g35593 not n20202 ; n20202_not
g35594 not n22101 ; n22101_not
g35595 not n15000 ; n15000_not
g35596 not n11103 ; n11103_not
g35597 not n21210 ; n21210_not
g35598 not n21021 ; n21021_not
g35599 not n10500 ; n10500_not
g35600 not n10122 ; n10122_not
g35601 not n11031 ; n11031_not
g35602 not n12111 ; n12111_not
g35603 not n10401 ; n10401_not
g35604 not n10113 ; n10113_not
g35605 not n11004 ; n11004_not
g35606 not n12210 ; n12210_not
g35607 not n12102 ; n12102_not
g35608 not n10104 ; n10104_not
g35609 not n24000 ; n24000_not
g35610 not n12201 ; n12201_not
g35611 not n20031 ; n20031_not
g35612 not n20040 ; n20040_not
g35613 not n12120 ; n12120_not
g35614 not n11022 ; n11022_not
g35615 not n11040 ; n11040_not
g35616 not n23010 ; n23010_not
g35617 not n13200 ; n13200_not
g35618 not n20301 ; n20301_not
g35619 not n11112 ; n11112_not
g35620 not n22200 ; n22200_not
g35621 not n11130 ; n11130_not
g35622 not n10131 ; n10131_not
g35623 not n20022 ; n20022_not
g35624 not n10140 ; n10140_not
g35625 not n13002 ; n13002_not
g35626 not n21040 ; n21040_not
g35627 not n12031 ; n12031_not
g35628 not n20131 ; n20131_not
g35629 not n12121 ; n12121_not
g35630 not n20122 ; n20122_not
g35631 not n20041 ; n20041_not
g35632 not n12400 ; n12400_not
g35633 not n22111 ; n22111_not
g35634 not n20113 ; n20113_not
g35635 not n12130 ; n12130_not
g35636 not n13111 ; n13111_not
g35637 not n10420 ; n10420_not
g35638 not n21013 ; n21013_not
g35639 not n10330 ; n10330_not
g35640 not n13120 ; n13120_not
g35641 not n24100 ; n24100_not
g35642 not n20050 ; n20050_not
g35643 not n13201 ; n13201_not
g35644 not n23020 ; n23020_not
g35645 not n10006 ; n10006_not
g35646 not n13210 ; n13210_not
g35647 not n10501 ; n10501_not
g35648 not n11500 ; n11500_not
g35649 not n21004 ; n21004_not
g35650 not n22120 ; n22120_not
g35651 not n20140 ; n20140_not
g35652 not n24010 ; n24010_not
g35653 not n13021 ; n13021_not
g35654 not n20032 ; n20032_not
g35655 not n12040 ; n12040_not
g35656 not n15010 ; n15010_not
g35657 not n10015 ; n10015_not
g35658 not n22003 ; n22003_not
g35659 not n13030 ; n13030_not
g35660 not n23110 ; n23110_not
g35661 not n12220 ; n12220_not
g35662 not n10321 ; n10321_not
g35663 not n10600 ; n10600_not
g35664 not n12013 ; n12013_not
g35665 not n10222 ; n10222_not
g35666 not n12310 ; n12310_not
g35667 not n20014 ; n20014_not
g35668 not n21022 ; n21022_not
g35669 not n21400 ; n21400_not
g35670 not n23200 ; n23200_not
g35671 not n12301 ; n12301_not
g35672 not n23002 ; n23002_not
g35673 not n12004 ; n12004_not
g35674 not n12022 ; n12022_not
g35675 not n12202 ; n12202_not
g35676 not n20005 ; n20005_not
g35677 not n10411 ; n10411_not
g35678 not n10510 ; n10510_not
g35679 not n21103 ; n21103_not
g35680 not n20104 ; n20104_not
g35681 not n10033 ; n10033_not
g35682 not n12112 ; n12112_not
g35683 not n10303 ; n10303_not
g35684 not n22021 ; n22021_not
g35685 not n13300 ; n13300_not
g35686 not n10402 ; n10402_not
g35687 not n13003 ; n13003_not
g35688 not n10312 ; n10312_not
g35689 not n12103 ; n12103_not
g35690 not n20311 ; n20311_not
g35691 not n14002 ; n14002_not
g35692 not n10114 ; n10114_not
g35693 not n15100 ; n15100_not
g35694 not n14200 ; n14200_not
g35695 not n16000 ; n16000_not
g35696 not n20230 ; n20230_not
g35697 not n11212 ; n11212_not
g35698 not n10051 ; n10051_not
g35699 not n11221 ; n11221_not
g35700 not n20320 ; n20320_not
g35701 not n11230 ; n11230_not
g35702 not n21310 ; n21310_not
g35703 not n11302 ; n11302_not
g35704 not n20221 ; n20221_not
g35705 not n11311 ; n11311_not
g35706 not n11320 ; n11320_not
g35707 not n10042 ; n10042_not
g35708 not n20203 ; n20203_not
g35709 not n10204 ; n10204_not
g35710 not n22210 ; n22210_not
g35711 not n11032 ; n11032_not
g35712 not n23011 ; n23011_not
g35713 not n11023 ; n11023_not
g35714 not n11041 ; n11041_not
g35715 not n24001 ; n24001_not
g35716 not n11014 ; n11014_not
g35717 not n10105 ; n10105_not
g35718 not n11005 ; n11005_not
g35719 not n11050 ; n11050_not
g35720 not n20302 ; n20302_not
g35721 not n21220 ; n21220_not
g35722 not n10123 ; n10123_not
g35723 not n21211 ; n21211_not
g35724 not n11104 ; n11104_not
g35725 not n11113 ; n11113_not
g35726 not n21202 ; n21202_not
g35727 not n11122 ; n11122_not
g35728 not n10141 ; n10141_not
g35729 not n10132 ; n10132_not
g35730 not n11131 ; n11131_not
g35731 not n10150 ; n10150_not
g35732 not n10240 ; n10240_not
g35733 not n14011 ; n14011_not
g35734 not n21121 ; n21121_not
g35735 not n14020 ; n14020_not
g35736 not n10231 ; n10231_not
g35737 not n20401 ; n20401_not
g35738 not n25000 ; n25000_not
g35739 not n11401 ; n11401_not
g35740 not n10213 ; n10213_not
g35741 not n14101 ; n14101_not
g35742 not n14110 ; n14110_not
g35743 not n10502 ; n10502_not
g35744 not n20204 ; n20204_not
g35745 not n11105 ; n11105_not
g35746 not n22130 ; n22130_not
g35747 not n11510 ; n11510_not
g35748 not n11024 ; n11024_not
g35749 not n20141 ; n20141_not
g35750 not n23021 ; n23021_not
g35751 not n14300 ; n14300_not
g35752 not n21023 ; n21023_not
g35753 not n12104 ; n12104_not
g35754 not n20303 ; n20303_not
g35755 not n11204 ; n11204_not
g35756 not n24110 ; n24110_not
g35757 not n23120 ; n23120_not
g35758 not n11231 ; n11231_not
g35759 not n22220 ; n22220_not
g35760 not n12050 ; n12050_not
g35761 not n20051 ; n20051_not
g35762 not n21005 ; n21005_not
g35763 not n13310 ; n13310_not
g35764 not n10520 ; n10520_not
g35765 not n11132 ; n11132_not
g35766 not n20501 ; n20501_not
g35767 not n11420 ; n11420_not
g35768 not n21014 ; n21014_not
g35769 not n22211 ; n22211_not
g35770 not n10511 ; n10511_not
g35771 not n24200 ; n24200_not
g35772 not n24011 ; n24011_not
g35773 not n14021 ; n14021_not
g35774 not n11222 ; n11222_not
g35775 not n22400 ; n22400_not
g35776 not n22310 ; n22310_not
g35777 not n12131 ; n12131_not
g35778 not n12140 ; n12140_not
g35779 not n23300 ; n23300_not
g35780 not n20420 ; n20420_not
g35781 not n20033 ; n20033_not
g35782 not n13220 ; n13220_not
g35783 not n10403 ; n10403_not
g35784 not n11033 ; n11033_not
g35785 not n20411 ; n20411_not
g35786 not n13211 ; n13211_not
g35787 not n13202 ; n13202_not
g35788 not n24002 ; n24002_not
g35789 not n12113 ; n12113_not
g35790 not n14012 ; n14012_not
g35791 not n14102 ; n14102_not
g35792 not n20042 ; n20042_not
g35793 not n13004 ; n13004_not
g35794 not n15110 ; n15110_not
g35795 not n11240 ; n11240_not
g35796 not n24101 ; n24101_not
g35797 not n12122 ; n12122_not
g35798 not n11015 ; n11015_not
g35799 not n23102 ; n23102_not
g35800 not n11042 ; n11042_not
g35801 not n20231 ; n20231_not
g35802 not n10610 ; n10610_not
g35803 not n11123 ; n11123_not
g35804 not n10601 ; n10601_not
g35805 not n10241 ; n10241_not
g35806 not n26000 ; n26000_not
g35807 not n11600 ; n11600_not
g35808 not n13103 ; n13103_not
g35809 not n20600 ; n20600_not
g35810 not n11060 ; n11060_not
g35811 not n20123 ; n20123_not
g35812 not n20240 ; n20240_not
g35813 not n13400 ; n13400_not
g35814 not n20213 ; n20213_not
g35815 not n23111 ; n23111_not
g35816 not n11312 ; n11312_not
g35817 not n22040 ; n22040_not
g35818 not n22022 ; n22022_not
g35819 not n11006 ; n11006_not
g35820 not n22112 ; n22112_not
g35821 not n11303 ; n11303_not
g35822 not n20024 ; n20024_not
g35823 not n23030 ; n23030_not
g35824 not n22013 ; n22013_not
g35825 not n22004 ; n22004_not
g35826 not n11321 ; n11321_not
g35827 not n14120 ; n14120_not
g35828 not n20330 ; n20330_not
g35829 not n14201 ; n14201_not
g35830 not n20312 ; n20312_not
g35831 not n14030 ; n14030_not
g35832 not n11150 ; n11150_not
g35833 not n12023 ; n12023_not
g35834 not n20510 ; n20510_not
g35835 not n12032 ; n12032_not
g35836 not n12041 ; n12041_not
g35837 not n11141 ; n11141_not
g35838 not n20114 ; n20114_not
g35839 not n16100 ; n16100_not
g35840 not n11213 ; n11213_not
g35841 not n10205 ; n10205_not
g35842 not n11411 ; n11411_not
g35843 not n20105 ; n20105_not
g35844 not n16001 ; n16001_not
g35845 not n24020 ; n24020_not
g35846 not n20132 ; n20132_not
g35847 not n12014 ; n12014_not
g35848 not n10133 ; n10133_not
g35849 not n12311 ; n12311_not
g35850 not n12410 ; n12410_not
g35851 not n21221 ; n21221_not
g35852 not n13022 ; n13022_not
g35853 not n21302 ; n21302_not
g35854 not n13130 ; n13130_not
g35855 not n21140 ; n21140_not
g35856 not n10070 ; n10070_not
g35857 not n21113 ; n21113_not
g35858 not n10106 ; n10106_not
g35859 not n10016 ; n10016_not
g35860 not n15011 ; n15011_not
g35861 not n12230 ; n12230_not
g35862 not n10142 ; n10142_not
g35863 not n10151 ; n10151_not
g35864 not n23012 ; n23012_not
g35865 not n12500 ; n12500_not
g35866 not n10322 ; n10322_not
g35867 not n10232 ; n10232_not
g35868 not n21203 ; n21203_not
g35869 not n21122 ; n21122_not
g35870 not n12401 ; n12401_not
g35871 not n12212 ; n12212_not
g35872 not n10124 ; n10124_not
g35873 not n10340 ; n10340_not
g35874 not n10025 ; n10025_not
g35875 not n17000 ; n17000_not
g35876 not n10304 ; n10304_not
g35877 not n12302 ; n12302_not
g35878 not n21212 ; n21212_not
g35879 not n23201 ; n23201_not
g35880 not n20015 ; n20015_not
g35881 not n10331 ; n10331_not
g35882 not n13112 ; n13112_not
g35883 not n15020 ; n15020_not
g35884 not n21311 ; n21311_not
g35885 not n10052 ; n10052_not
g35886 not n21320 ; n21320_not
g35887 not n10061 ; n10061_not
g35888 not n10115 ; n10115_not
g35889 not n23003 ; n23003_not
g35890 not n10250 ; n10250_not
g35891 not n21410 ; n21410_not
g35892 not n21401 ; n21401_not
g35893 not n10007 ; n10007_not
g35894 not n21032 ; n21032_not
g35895 not n21041 ; n21041_not
g35896 not n13040 ; n13040_not
g35897 not n10214 ; n10214_not
g35898 not n10313 ; n10313_not
g35899 not n21500 ; n21500_not
g35900 not n25010 ; n25010_not
g35901 not n10430 ; n10430_not
g35902 not n25001 ; n25001_not
g35903 not n21104 ; n21104_not
g35904 not n10160 ; n10160_not
g35905 not n13031 ; n13031_not
g35906 not n20006 ; n20006_not
g35907 not n10034 ; n10034_not
g35908 not n10412 ; n10412_not
g35909 not n10043 ; n10043_not
g35910 not n21131 ; n21131_not
g35911 not n25100 ; n25100_not
g35912 not n21230 ; n21230_not
g35913 not n15101 ; n15101_not
g35914 not n10223 ; n10223_not
g35915 not n20250 ; n20250_not
g35916 not n20502 ; n20502_not
g35917 not n10710 ; n10710_not
g35918 not n12411 ; n12411_not
g35919 not n20106 ; n20106_not
g35920 not n11160 ; n11160_not
g35921 not n25110 ; n25110_not
g35922 not n26100 ; n26100_not
g35923 not n15021 ; n15021_not
g35924 not n20304 ; n20304_not
g35925 not n20313 ; n20313_not
g35926 not n10260 ; n10260_not
g35927 not n24201 ; n24201_not
g35928 not n20142 ; n20142_not
g35929 not n11700 ; n11700_not
g35930 not n14202 ; n14202_not
g35931 not n12303 ; n12303_not
g35932 not n12240 ; n12240_not
g35933 not n15012 ; n15012_not
g35934 not n22500 ; n22500_not
g35935 not n16002 ; n16002_not
g35936 not n20520 ; n20520_not
g35937 not n10053 ; n10053_not
g35938 not n15300 ; n15300_not
g35939 not n11610 ; n11610_not
g35940 not n13032 ; n13032_not
g35941 not n18000 ; n18000_not
g35942 not n20124 ; n20124_not
g35943 not n12402 ; n12402_not
g35944 not n25101 ; n25101_not
g35945 not n22311 ; n22311_not
g35946 not n11601 ; n11601_not
g35947 not n21411 ; n21411_not
g35948 not n11205 ; n11205_not
g35949 not n24210 ; n24210_not
g35950 not n17001 ; n17001_not
g35951 not n24012 ; n24012_not
g35952 not n21105 ; n21105_not
g35953 not n22221 ; n22221_not
g35954 not n14220 ; n14220_not
g35955 not n10341 ; n10341_not
g35956 not n22113 ; n22113_not
g35957 not n23103 ; n23103_not
g35958 not n22104 ; n22104_not
g35959 not n15003 ; n15003_not
g35960 not n13041 ; n13041_not
g35961 not n14103 ; n14103_not
g35962 not n25011 ; n25011_not
g35963 not n21330 ; n21330_not
g35964 not n10215 ; n10215_not
g35965 not n11106 ; n11106_not
g35966 not n20331 ; n20331_not
g35967 not n21132 ; n21132_not
g35968 not n14040 ; n14040_not
g35969 not n25002 ; n25002_not
g35970 not n20232 ; n20232_not
g35971 not n11412 ; n11412_not
g35972 not n10224 ; n10224_not
g35973 not n20340 ; n20340_not
g35974 not n14031 ; n14031_not
g35975 not n21123 ; n21123_not
g35976 not n20403 ; n20403_not
g35977 not n11052 ; n11052_not
g35978 not n11421 ; n11421_not
g35979 not n10440 ; n10440_not
g35980 not n10233 ; n10233_not
g35981 not n23040 ; n23040_not
g35982 not n22302 ; n22302_not
g35983 not n11304 ; n11304_not
g35984 not n20214 ; n20214_not
g35985 not n21150 ; n21150_not
g35986 not n20223 ; n20223_not
g35987 not n25020 ; n25020_not
g35988 not n11322 ; n11322_not
g35989 not n20205 ; n20205_not
g35990 not n10044 ; n10044_not
g35991 not n11313 ; n11313_not
g35992 not n12510 ; n12510_not
g35993 not n11331 ; n11331_not
g35994 not n10206 ; n10206_not
g35995 not n23112 ; n23112_not
g35996 not n11340 ; n11340_not
g35997 not n22005 ; n22005_not
g35998 not n14121 ; n14121_not
g35999 not n22320 ; n22320_not
g36000 not n11232 ; n11232_not
g36001 not n22410 ; n22410_not
g36002 not n20160 ; n20160_not
g36003 not n14400 ; n14400_not
g36004 not n21114 ; n21114_not
g36005 not n21312 ; n21312_not
g36006 not n13014 ; n13014_not
g36007 not n22212 ; n22212_not
g36008 not n11511 ; n11511_not
g36009 not n21024 ; n21024_not
g36010 not n20430 ; n20430_not
g36011 not n11520 ; n11520_not
g36012 not n24120 ; n24120_not
g36013 not n11223 ; n11223_not
g36014 not n16200 ; n16200_not
g36015 not n21303 ; n21303_not
g36016 not n16101 ; n16101_not
g36017 not n12420 ; n12420_not
g36018 not n22131 ; n22131_not
g36019 not n10170 ; n10170_not
g36020 not n22230 ; n22230_not
g36021 not n11250 ; n11250_not
g36022 not n11430 ; n11430_not
g36023 not n21321 ; n21321_not
g36024 not n11241 ; n11241_not
g36025 not n14013 ; n14013_not
g36026 not n21141 ; n21141_not
g36027 not n15030 ; n15030_not
g36028 not n10017 ; n10017_not
g36029 not n14004 ; n14004_not
g36030 not n21402 ; n21402_not
g36031 not n20412 ; n20412_not
g36032 not n20421 ; n20421_not
g36033 not n13005 ; n13005_not
g36034 not n16110 ; n16110_not
g36035 not n10251 ; n10251_not
g36036 not n24102 ; n24102_not
g36037 not n11043 ; n11043_not
g36038 not n12033 ; n12033_not
g36039 not n13113 ; n13113_not
g36040 not n12042 ; n12042_not
g36041 not n21060 ; n21060_not
g36042 not n13320 ; n13320_not
g36043 not n23130 ; n23130_not
g36044 not n24003 ; n24003_not
g36045 not n12051 ; n12051_not
g36046 not n10116 ; n10116_not
g36047 not n20052 ; n20052_not
g36048 not n23310 ; n23310_not
g36049 not n10530 ; n10530_not
g36050 not n21051 ; n21051_not
g36051 not n12114 ; n12114_not
g36052 not n21006 ; n21006_not
g36053 not n23022 ; n23022_not
g36054 not n13311 ; n13311_not
g36055 not n12132 ; n12132_not
g36056 not n13302 ; n13302_not
g36057 not n20070 ; n20070_not
g36058 not n10431 ; n10431_not
g36059 not n20034 ; n20034_not
g36060 not n23400 ; n23400_not
g36061 not n10350 ; n10350_not
g36062 not n10062 ; n10062_not
g36063 not n12015 ; n12015_not
g36064 not n12141 ; n12141_not
g36065 not n23202 ; n23202_not
g36066 not n20016 ; n20016_not
g36067 not n21213 ; n21213_not
g36068 not n11070 ; n11070_not
g36069 not n21231 ; n21231_not
g36070 not n11061 ; n11061_not
g36071 not n23301 ; n23301_not
g36072 not n21501 ; n21501_not
g36073 not n12231 ; n12231_not
g36074 not n21042 ; n21042_not
g36075 not n12213 ; n12213_not
g36076 not n27000 ; n27000_not
g36077 not n23031 ; n23031_not
g36078 not n23013 ; n23013_not
g36079 not n12123 ; n12123_not
g36080 not n11016 ; n11016_not
g36081 not n12105 ; n12105_not
g36082 not n15210 ; n15210_not
g36083 not n10404 ; n10404_not
g36084 not n20043 ; n20043_not
g36085 not n10413 ; n10413_not
g36086 not n12060 ; n12060_not
g36087 not n10521 ; n10521_not
g36088 not n23121 ; n23121_not
g36089 not n10422 ; n10422_not
g36090 not n23220 ; n23220_not
g36091 not n21015 ; n21015_not
g36092 not n13131 ; n13131_not
g36093 not n21222 ; n21222_not
g36094 not n21600 ; n21600_not
g36095 not n11007 ; n11007_not
g36096 not n20025 ; n20025_not
g36097 not n11034 ; n11034_not
g36098 not n10503 ; n10503_not
g36099 not n13212 ; n13212_not
g36100 not n12600 ; n12600_not
g36101 not n15120 ; n15120_not
g36102 not n10125 ; n10125_not
g36103 not n11133 ; n11133_not
g36104 not n10314 ; n10314_not
g36105 not n10305 ; n10305_not
g36106 not n10611 ; n10611_not
g36107 not n10026 ; n10026_not
g36108 not n20610 ; n20610_not
g36109 not n23004 ; n23004_not
g36110 not n20601 ; n20601_not
g36111 not n10602 ; n10602_not
g36112 not n13410 ; n13410_not
g36113 not n22023 ; n22023_not
g36114 not n11142 ; n11142_not
g36115 not n10080 ; n10080_not
g36116 not n22032 ; n22032_not
g36117 not n22014 ; n22014_not
g36118 not n13221 ; n13221_not
g36119 not n10152 ; n10152_not
g36120 not n15111 ; n15111_not
g36121 not n15102 ; n15102_not
g36122 not n21510 ; n21510_not
g36123 not n10620 ; n10620_not
g36124 not n21033 ; n21033_not
g36125 not n13500 ; n13500_not
g36126 not n10134 ; n10134_not
g36127 not n22203 ; n22203_not
g36128 not n10323 ; n10323_not
g36129 not n25200 ; n25200_not
g36130 not n21240 ; n21240_not
g36131 not n12330 ; n12330_not
g36132 not n14310 ; n14310_not
g36133 not n21204 ; n21204_not
g36134 not n10332 ; n10332_not
g36135 not n13203 ; n13203_not
g36136 not n13401 ; n13401_not
g36137 not n13104 ; n13104_not
g36138 not n20700 ; n20700_not
g36139 not n10143 ; n10143_not
g36140 not n26010 ; n26010_not
g36141 not n22041 ; n22041_not
g36142 not n11124 ; n11124_not
g36143 not n11025 ; n11025_not
g36144 not n12312 ; n12312_not
g36145 not n12150 ; n12150_not
g36146 not n13230 ; n13230_not
g36147 not n14301 ; n14301_not
g36148 not n10900 ; n10900_not
g36149 not n21340 ; n21340_not
g36150 not n11305 ; n11305_not
g36151 not n17110 ; n17110_not
g36152 not n12700 ; n12700_not
g36153 not n17101 ; n17101_not
g36154 not n25030 ; n25030_not
g36155 not n21250 ; n21250_not
g36156 not n12511 ; n12511_not
g36157 not n21232 ; n21232_not
g36158 not n14122 ; n14122_not
g36159 not n21331 ; n21331_not
g36160 not n21043 ; n21043_not
g36161 not n11035 ; n11035_not
g36162 not n11044 ; n11044_not
g36163 not n12502 ; n12502_not
g36164 not n20332 ; n20332_not
g36165 not n25201 ; n25201_not
g36166 not n14131 ; n14131_not
g36167 not n21322 ; n21322_not
g36168 not n12403 ; n12403_not
g36169 not n12520 ; n12520_not
g36170 not n23023 ; n23023_not
g36171 not n25120 ; n25120_not
g36172 not n21205 ; n21205_not
g36173 not n14230 ; n14230_not
g36174 not n11206 ; n11206_not
g36175 not n11116 ; n11116_not
g36176 not n12610 ; n12610_not
g36177 not n11125 ; n11125_not
g36178 not n15301 ; n15301_not
g36179 not n12601 ; n12601_not
g36180 not n17020 ; n17020_not
g36181 not n20314 ; n20314_not
g36182 not n18001 ; n18001_not
g36183 not n24022 ; n24022_not
g36184 not n20305 ; n20305_not
g36185 not n18010 ; n18010_not
g36186 not n24013 ; n24013_not
g36187 not n11143 ; n11143_not
g36188 not n17002 ; n17002_not
g36189 not n17200 ; n17200_not
g36190 not n25111 ; n25111_not
g36191 not n14203 ; n14203_not
g36192 not n14104 ; n14104_not
g36193 not n14212 ; n14212_not
g36194 not n25300 ; n25300_not
g36195 not n11161 ; n11161_not
g36196 not n14140 ; n14140_not
g36197 not n16120 ; n16120_not
g36198 not n11260 ; n11260_not
g36199 not n11251 ; n11251_not
g36200 not n21214 ; n21214_not
g36201 not n21223 ; n21223_not
g36202 not n20323 ; n20323_not
g36203 not n24040 ; n24040_not
g36204 not n11134 ; n11134_not
g36205 not n11242 ; n11242_not
g36206 not n11053 ; n11053_not
g36207 not n16111 ; n16111_not
g36208 not n11233 ; n11233_not
g36209 not n22150 ; n22150_not
g36210 not n11170 ; n11170_not
g36211 not n16102 ; n16102_not
g36212 not n24004 ; n24004_not
g36213 not n11062 ; n11062_not
g36214 not n11224 ; n11224_not
g36215 not n21304 ; n21304_not
g36216 not n12241 ; n12241_not
g36217 not n11080 ; n11080_not
g36218 not n24031 ; n24031_not
g36219 not n22204 ; n22204_not
g36220 not n20341 ; n20341_not
g36221 not n20800 ; n20800_not
g36222 not n11530 ; n11530_not
g36223 not n13510 ; n13510_not
g36224 not n13501 ; n13501_not
g36225 not n13114 ; n13114_not
g36226 not n13132 ; n13132_not
g36227 not n13240 ; n13240_not
g36228 not n13420 ; n13420_not
g36229 not n21700 ; n21700_not
g36230 not n13411 ; n13411_not
g36231 not n13402 ; n13402_not
g36232 not n24400 ; n24400_not
g36233 not n20701 ; n20701_not
g36234 not n13105 ; n13105_not
g36235 not n12007 ; n12007_not
g36236 not n23032 ; n23032_not
g36237 not n21070 ; n21070_not
g36238 not n12016 ; n12016_not
g36239 not n21610 ; n21610_not
g36240 not n22042 ; n22042_not
g36241 not n12331 ; n12331_not
g36242 not n20602 ; n20602_not
g36243 not n22033 ; n22033_not
g36244 not n20611 ; n20611_not
g36245 not n22024 ; n22024_not
g36246 not n13042 ; n13042_not
g36247 not n12322 ; n12322_not
g36248 not n22015 ; n22015_not
g36249 not n20422 ; n20422_not
g36250 not n15202 ; n15202_not
g36251 not n26020 ; n26020_not
g36252 not n11800 ; n11800_not
g36253 not n22006 ; n22006_not
g36254 not n11422 ; n11422_not
g36255 not n27100 ; n27100_not
g36256 not n12313 ; n12313_not
g36257 not n26011 ; n26011_not
g36258 not n13600 ; n13600_not
g36259 not n26002 ; n26002_not
g36260 not n12214 ; n12214_not
g36261 not n12205 ; n12205_not
g36262 not n12115 ; n12115_not
g36263 not n12133 ; n12133_not
g36264 not n21520 ; n21520_not
g36265 not n21502 ; n21502_not
g36266 not n21511 ; n21511_not
g36267 not n12142 ; n12142_not
g36268 not n21025 ; n21025_not
g36269 not n13231 ; n13231_not
g36270 not n12151 ; n12151_not
g36271 not n13222 ; n13222_not
g36272 not n15211 ; n15211_not
g36273 not n12160 ; n12160_not
g36274 not n15310 ; n15310_not
g36275 not n21034 ; n21034_not
g36276 not n13006 ; n13006_not
g36277 not n21061 ; n21061_not
g36278 not n12052 ; n12052_not
g36279 not n13321 ; n13321_not
g36280 not n13123 ; n13123_not
g36281 not n21007 ; n21007_not
g36282 not n21052 ; n21052_not
g36283 not n12061 ; n12061_not
g36284 not n12070 ; n12070_not
g36285 not n13303 ; n13303_not
g36286 not n12250 ; n12250_not
g36287 not n21601 ; n21601_not
g36288 not n13141 ; n13141_not
g36289 not n12232 ; n12232_not
g36290 not n13150 ; n13150_not
g36291 not n12223 ; n12223_not
g36292 not n21124 ; n21124_not
g36293 not n11404 ; n11404_not
g36294 not n11413 ; n11413_not
g36295 not n14032 ; n14032_not
g36296 not n14023 ; n14023_not
g36297 not n11431 ; n11431_not
g36298 not n20404 ; n20404_not
g36299 not n23104 ; n23104_not
g36300 not n11440 ; n11440_not
g36301 not n14014 ; n14014_not
g36302 not n14005 ; n14005_not
g36303 not n20413 ; n20413_not
g36304 not n26200 ; n26200_not
g36305 not n21403 ; n21403_not
g36306 not n12430 ; n12430_not
g36307 not n21115 ; n21115_not
g36308 not n24103 ; n24103_not
g36309 not n20431 ; n20431_not
g36310 not n21142 ; n21142_not
g36311 not n21151 ; n21151_not
g36312 not n11314 ; n11314_not
g36313 not n25021 ; n25021_not
g36314 not n25012 ; n25012_not
g36315 not n11323 ; n11323_not
g36316 not n14113 ; n14113_not
g36317 not n21133 ; n21133_not
g36318 not n11332 ; n11332_not
g36319 not n20044 ; n20044_not
g36320 not n11341 ; n11341_not
g36321 not n11350 ; n11350_not
g36322 not n20350 ; n20350_not
g36323 not n11107 ; n11107_not
g36324 not n14041 ; n14041_not
g36325 not n11071 ; n11071_not
g36326 not n14050 ; n14050_not
g36327 not n25003 ; n25003_not
g36328 not n20521 ; n20521_not
g36329 not n11611 ; n11611_not
g36330 not n12340 ; n12340_not
g36331 not n21412 ; n21412_not
g36332 not n13033 ; n13033_not
g36333 not n11620 ; n11620_not
g36334 not n22105 ; n22105_not
g36335 not n21421 ; n21421_not
g36336 not n21106 ; n21106_not
g36337 not n20530 ; n20530_not
g36338 not n16300 ; n16300_not
g36339 not n20242 ; n20242_not
g36340 not n26101 ; n26101_not
g36341 not n24310 ; n24310_not
g36342 not n11701 ; n11701_not
g36343 not n22060 ; n22060_not
g36344 not n11710 ; n11710_not
g36345 not n13060 ; n13060_not
g36346 not n22051 ; n22051_not
g36347 not n21430 ; n21430_not
g36348 not n13015 ; n13015_not
g36349 not n11503 ; n11503_not
g36350 not n20440 ; n20440_not
g36351 not n11512 ; n11512_not
g36352 not n22141 ; n22141_not
g36353 not n24121 ; n24121_not
g36354 not n16201 ; n16201_not
g36355 not n16210 ; n16210_not
g36356 not n11521 ; n11521_not
g36357 not n12421 ; n12421_not
g36358 not n22132 ; n22132_not
g36359 not n22123 ; n22123_not
g36360 not n12412 ; n12412_not
g36361 not n12304 ; n12304_not
g36362 not n22114 ; n22114_not
g36363 not n24211 ; n24211_not
g36364 not n20512 ; n20512_not
g36365 not n11602 ; n11602_not
g36366 not n24220 ; n24220_not
g36367 not n15400 ; n15400_not
g36368 not n23140 ; n23140_not
g36369 not n14221 ; n14221_not
g36370 not n20224 ; n20224_not
g36371 not n10540 ; n10540_not
g36372 not n20215 ; n20215_not
g36373 not n19000 ; n19000_not
g36374 not n20206 ; n20206_not
g36375 not n22303 ; n22303_not
g36376 not n10054 ; n10054_not
g36377 not n23041 ; n23041_not
g36378 not n22312 ; n22312_not
g36379 not n22321 ; n22321_not
g36380 not n20053 ; n20053_not
g36381 not n10045 ; n10045_not
g36382 not n10216 ; n10216_not
g36383 not n15040 ; n15040_not
g36384 not n10018 ; n10018_not
g36385 not n10234 ; n10234_not
g36386 not n10225 ; n10225_not
g36387 not n10522 ; n10522_not
g36388 not n22600 ; n22600_not
g36389 not n10243 ; n10243_not
g36390 not n15031 ; n15031_not
g36391 not n10252 ; n10252_not
g36392 not n10810 ; n10810_not
g36393 not n15022 ; n15022_not
g36394 not n10801 ; n10801_not
g36395 not n10270 ; n10270_not
g36396 not n10261 ; n10261_not
g36397 not n10063 ; n10063_not
g36398 not n23131 ; n23131_not
g36399 not n10126 ; n10126_not
g36400 not n20251 ; n20251_not
g36401 not n10135 ; n10135_not
g36402 not n16012 ; n16012_not
g36403 not n10144 ; n10144_not
g36404 not n15103 ; n15103_not
g36405 not n16003 ; n16003_not
g36406 not n23014 ; n23014_not
g36407 not n22222 ; n22222_not
g36408 not n22231 ; n22231_not
g36409 not n14410 ; n14410_not
g36410 not n10180 ; n10180_not
g36411 not n20062 ; n20062_not
g36412 not n20233 ; n20233_not
g36413 not n10171 ; n10171_not
g36414 not n10090 ; n10090_not
g36415 not n23401 ; n23401_not
g36416 not n23203 ; n23203_not
g36417 not n14401 ; n14401_not
g36418 not n10162 ; n10162_not
g36419 not n20017 ; n20017_not
g36420 not n22402 ; n22402_not
g36421 not n23500 ; n23500_not
g36422 not n23320 ; n23320_not
g36423 not n10621 ; n10621_not
g36424 not n20125 ; n20125_not
g36425 not n23212 ; n23212_not
g36426 not n10630 ; n10630_not
g36427 not n22501 ; n22501_not
g36428 not n23221 ; n23221_not
g36429 not n20107 ; n20107_not
g36430 not n23230 ; n23230_not
g36431 not n23311 ; n23311_not
g36432 not n10342 ; n10342_not
g36433 not n23302 ; n23302_not
g36434 not n10414 ; n10414_not
g36435 not n10423 ; n10423_not
g36436 not n22510 ; n22510_not
g36437 not n20026 ; n20026_not
g36438 not n10432 ; n10432_not
g36439 not n10405 ; n10405_not
g36440 not n27010 ; n27010_not
g36441 not n10441 ; n10441_not
g36442 not n10450 ; n10450_not
g36443 not n15004 ; n15004_not
g36444 not n20161 ; n20161_not
g36445 not n22240 ; n22240_not
g36446 not n22411 ; n22411_not
g36447 not n10603 ; n10603_not
g36448 not n10504 ; n10504_not
g36449 not n22420 ; n22420_not
g36450 not n23113 ; n23113_not
g36451 not n20152 ; n20152_not
g36452 not n23410 ; n23410_not
g36453 not n27001 ; n27001_not
g36454 not n10612 ; n10612_not
g36455 not n10351 ; n10351_not
g36456 not n10702 ; n10702_not
g36457 not n10333 ; n10333_not
g36458 not n10711 ; n10711_not
g36459 not n20143 ; n20143_not
g36460 not n10720 ; n10720_not
g36461 not n10324 ; n10324_not
g36462 not n10027 ; n10027_not
g36463 not n10315 ; n10315_not
g36464 not n10306 ; n10306_not
g36465 not n18100 ; n18100_not
g36466 not n10117 ; n10117_not
g36467 not n16021 ; n16021_not
g36468 not n11008 ; n11008_not
g36469 not n14320 ; n14320_not
g36470 not n10081 ; n10081_not
g36471 not n11017 ; n11017_not
g36472 not n20260 ; n20260_not
g36473 not n22213 ; n22213_not
g36474 not n14311 ; n14311_not
g36475 not n15121 ; n15121_not
g36476 not n20071 ; n20071_not
g36477 not n14302 ; n14302_not
g36478 not n23005 ; n23005_not
g36479 not n15112 ; n15112_not
g36480 not n12341 ; n12341_not
g36481 not n15230 ; n15230_not
g36482 not n21440 ; n21440_not
g36483 not n10730 ; n10730_not
g36484 not n22430 ; n22430_not
g36485 not n16211 ; n16211_not
g36486 not n25013 ; n25013_not
g36487 not n20315 ; n20315_not
g36488 not n27002 ; n27002_not
g36489 not n11540 ; n11540_not
g36490 not n11522 ; n11522_not
g36491 not n13043 ; n13043_not
g36492 not n24140 ; n24140_not
g36493 not n11027 ; n11027_not
g36494 not n22421 ; n22421_not
g36495 not n11801 ; n11801_not
g36496 not n11513 ; n11513_not
g36497 not n10451 ; n10451_not
g36498 not n13061 ; n13061_not
g36499 not n13070 ; n13070_not
g36500 not n15302 ; n15302_not
g36501 not n20009 ; n20009_not
g36502 not n20441 ; n20441_not
g36503 not n23042 ; n23042_not
g36504 not n20153 ; n20153_not
g36505 not n11810 ; n11810_not
g36506 not n24122 ; n24122_not
g36507 not n12350 ; n12350_not
g36508 not n15203 ; n15203_not
g36509 not n21431 ; n21431_not
g36510 not n12620 ; n12620_not
g36511 not n16202 ; n16202_not
g36512 not n11342 ; n11342_not
g36513 not n23105 ; n23105_not
g36514 not n21026 ; n21026_not
g36515 not n12314 ; n12314_not
g36516 not n25202 ; n25202_not
g36517 not n21701 ; n21701_not
g36518 not n10325 ; n10325_not
g36519 not n22124 ; n22124_not
g36520 not n23015 ; n23015_not
g36521 not n24041 ; n24041_not
g36522 not n20045 ; n20045_not
g36523 not n15122 ; n15122_not
g36524 not n20144 ; n20144_not
g36525 not n11063 ; n11063_not
g36526 not n24203 ; n24203_not
g36527 not n12305 ; n12305_not
g36528 not n10712 ; n10712_not
g36529 not n20072 ; n20072_not
g36530 not n10028 ; n10028_not
g36531 not n24005 ; n24005_not
g36532 not n10307 ; n10307_not
g36533 not n20603 ; n20603_not
g36534 not n10613 ; n10613_not
g36535 not n16220 ; n16220_not
g36536 not n12323 ; n12323_not
g36537 not n22133 ; n22133_not
g36538 not n23600 ; n23600_not
g36539 not n16040 ; n16040_not
g36540 not n14600 ; n14600_not
g36541 not n25040 ; n25040_not
g36542 not n10316 ; n10316_not
g36543 not n11225 ; n11225_not
g36544 not n21080 ; n21080_not
g36545 not n10280 ; n10280_not
g36546 not n11450 ; n11450_not
g36547 not n15320 ; n15320_not
g36548 not n10514 ; n10514_not
g36549 not n17300 ; n17300_not
g36550 not n20702 ; n20702_not
g36551 not n23330 ; n23330_not
g36552 not n21107 ; n21107_not
g36553 not n14006 ; n14006_not
g36554 not n14150 ; n14150_not
g36555 not n12080 ; n12080_not
g36556 not n26012 ; n26012_not
g36557 not n10460 ; n10460_not
g36558 not n20171 ; n20171_not
g36559 not n26201 ; n26201_not
g36560 not n15005 ; n15005_not
g36561 not n22205 ; n22205_not
g36562 not n22151 ; n22151_not
g36563 not n10622 ; n10622_not
g36564 not n10271 ; n10271_not
g36565 not n11090 ; n11090_not
g36566 not n12071 ; n12071_not
g36567 not n11432 ; n11432_not
g36568 not n13610 ; n13610_not
g36569 not n19001 ; n19001_not
g36570 not n14510 ; n14510_not
g36571 not n12404 ; n12404_not
g36572 not n14204 ; n14204_not
g36573 not n11441 ; n11441_not
g36574 not n14015 ; n14015_not
g36575 not n20405 ; n20405_not
g36576 not n14141 ; n14141_not
g36577 not n13025 ; n13025_not
g36578 not n18101 ; n18101_not
g36579 not n22142 ; n22142_not
g36580 not n10505 ; n10505_not
g36581 not n20432 ; n20432_not
g36582 not n14303 ; n14303_not
g36583 not n21602 ; n21602_not
g36584 not n11207 ; n11207_not
g36585 not n20306 ; n20306_not
g36586 not n24113 ; n24113_not
g36587 not n24410 ; n24410_not
g36588 not n21233 ; n21233_not
g36589 not n11504 ; n11504_not
g36590 not n21422 ; n21422_not
g36591 not n23051 ; n23051_not
g36592 not n15221 ; n15221_not
g36593 not n13034 ; n13034_not
g36594 not n22034 ; n22034_not
g36595 not n22403 ; n22403_not
g36596 not n21413 ; n21413_not
g36597 not n20162 ; n20162_not
g36598 not n27110 ; n27110_not
g36599 not n23060 ; n23060_not
g36600 not n13223 ; n13223_not
g36601 not n17102 ; n17102_not
g36602 not n11081 ; n11081_not
g36603 not n20423 ; n20423_not
g36604 not n10037 ; n10037_not
g36605 not n24104 ; n24104_not
g36606 not n13052 ; n13052_not
g36607 not n13160 ; n13160_not
g36608 not n12134 ; n12134_not
g36609 not n12215 ; n12215_not
g36610 not n21521 ; n21521_not
g36611 not n27020 ; n27020_not
g36612 not n23240 ; n23240_not
g36613 not n15140 ; n15140_not
g36614 not n20630 ; n20630_not
g36615 not n13412 ; n13412_not
g36616 not n24302 ; n24302_not
g36617 not n20900 ; n20900_not
g36618 not n10631 ; n10631_not
g36619 not n26102 ; n26102_not
g36620 not n12206 ; n12206_not
g36621 not n21044 ; n21044_not
g36622 not n10406 ; n10406_not
g36623 not n13250 ; n13250_not
g36624 not n13142 ; n13142_not
g36625 not n20612 ; n20612_not
g36626 not n16301 ; n16301_not
g36627 not n23312 ; n23312_not
g36628 not n13007 ; n13007_not
g36629 not n22502 ; n22502_not
g36630 not n27011 ; n27011_not
g36631 not n13151 ; n13151_not
g36632 not n12170 ; n12170_not
g36633 not n12224 ; n12224_not
g36634 not n22052 ; n22052_not
g36635 not n16310 ; n16310_not
g36636 not n15041 ; n15041_not
g36637 not n10433 ; n10433_not
g36638 not n22025 ; n22025_not
g36639 not n10442 ; n10442_not
g36640 not n13700 ; n13700_not
g36641 not n11711 ; n11711_not
g36642 not n23510 ; n23510_not
g36643 not n24320 ; n24320_not
g36644 not n20027 ; n20027_not
g36645 not n13205 ; n13205_not
g36646 not n11720 ; n11720_not
g36647 not n12143 ; n12143_not
g36648 not n23411 ; n23411_not
g36649 not n12701 ; n12701_not
g36650 not n23114 ; n23114_not
g36651 not n10415 ; n10415_not
g36652 not n12710 ; n12710_not
g36653 not n10424 ; n10424_not
g36654 not n24311 ; n24311_not
g36655 not n13241 ; n13241_not
g36656 not n22061 ; n22061_not
g36657 not n15212 ; n15212_not
g36658 not n22214 ; n22214_not
g36659 not n16400 ; n16400_not
g36660 not n23303 ; n23303_not
g36661 not n11702 ; n11702_not
g36662 not n21503 ; n21503_not
g36663 not n17120 ; n17120_not
g36664 not n21512 ; n21512_not
g36665 not n11036 ; n11036_not
g36666 not n21062 ; n21062_not
g36667 not n24230 ; n24230_not
g36668 not n11603 ; n11603_not
g36669 not n20135 ; n20135_not
g36670 not n23204 ; n23204_not
g36671 not n10640 ; n10640_not
g36672 not n20522 ; n20522_not
g36673 not n20126 ; n20126_not
g36674 not n11612 ; n11612_not
g36675 not n24221 ; n24221_not
g36676 not n23213 ; n23213_not
g36677 not n12116 ; n12116_not
g36678 not n24401 ; n24401_not
g36679 not n20018 ; n20018_not
g36680 not n20081 ; n20081_not
g36681 not n20504 ; n20504_not
g36682 not n13106 ; n13106_not
g36683 not n10343 ; n10343_not
g36684 not n10082 ; n10082_not
g36685 not n22115 ; n22115_not
g36686 not n17111 ; n17111_not
g36687 not n10703 ; n10703_not
g36688 not n21071 ; n21071_not
g36689 not n10352 ; n10352_not
g36690 not n12161 ; n12161_not
g36691 not n24212 ; n24212_not
g36692 not n11234 ; n11234_not
g36693 not n11054 ; n11054_not
g36694 not n20117 ; n20117_not
g36695 not n11009 ; n11009_not
g36696 not n12260 ; n12260_not
g36697 not n20108 ; n20108_not
g36698 not n12251 ; n12251_not
g36699 not n10154 ; n10154_not
g36700 not n15104 ; n15104_not
g36701 not n11018 ; n11018_not
g36702 not n23222 ; n23222_not
g36703 not n13133 ; n13133_not
g36704 not n12242 ; n12242_not
g36705 not n21530 ; n21530_not
g36706 not n12152 ; n12152_not
g36707 not n11045 ; n11045_not
g36708 not n25220 ; n25220_not
g36709 not n13115 ; n13115_not
g36710 not n23501 ; n23501_not
g36711 not n10370 ; n10370_not
g36712 not n13124 ; n13124_not
g36713 not n11621 ; n11621_not
g36714 not n21053 ; n21053_not
g36715 not n22520 ; n22520_not
g36716 not n20513 ; n20513_not
g36717 not n11630 ; n11630_not
g36718 not n22043 ; n22043_not
g36719 not n25400 ; n25400_not
g36720 not n23420 ; n23420_not
g36721 not n22016 ; n22016_not
g36722 not n22106 ; n22106_not
g36723 not n14411 ; n14411_not
g36724 not n11261 ; n11261_not
g36725 not n12026 ; n12026_not
g36726 not n22610 ; n22610_not
g36727 not n20324 ; n20324_not
g36728 not n20234 ; n20234_not
g36729 not n10109 ; n10109_not
g36730 not n16121 ; n16121_not
g36731 not n13331 ; n13331_not
g36732 not n11270 ; n11270_not
g36733 not n20090 ; n20090_not
g36734 not n14420 ; n14420_not
g36735 not n13511 ; n13511_not
g36736 not n21611 ; n21611_not
g36737 not n10091 ; n10091_not
g36738 not n14402 ; n14402_not
g36739 not n17210 ; n17210_not
g36740 not n10163 ; n10163_not
g36741 not n14222 ; n14222_not
g36742 not n11135 ; n11135_not
g36743 not n11243 ; n11243_not
g36744 not n10172 ; n10172_not
g36745 not n20063 ; n20063_not
g36746 not n13502 ; n13502_not
g36747 not n12017 ; n12017_not
g36748 not n11126 ; n11126_not
g36749 not n20261 ; n20261_not
g36750 not n23141 ; n23141_not
g36751 not n21305 ; n21305_not
g36752 not n11252 ; n11252_not
g36753 not n10541 ; n10541_not
g36754 not n25022 ; n25022_not
g36755 not n12035 ; n12035_not
g36756 not n20225 ; n20225_not
g36757 not n21224 ; n21224_not
g36758 not n20207 ; n20207_not
g36759 not n11306 ; n11306_not
g36760 not n25031 ; n25031_not
g36761 not n14114 ; n14114_not
g36762 not n12512 ; n12512_not
g36763 not n14330 ; n14330_not
g36764 not n20216 ; n20216_not
g36765 not n11315 ; n11315_not
g36766 not n10055 ; n10055_not
g36767 not n14312 ; n14312_not
g36768 not n13520 ; n13520_not
g36769 not n10073 ; n10073_not
g36770 not n17030 ; n17030_not
g36771 not n12530 ; n12530_not
g36772 not n11117 ; n11117_not
g36773 not n24050 ; n24050_not
g36774 not n21323 ; n21323_not
g36775 not n14123 ; n14123_not
g36776 not n25130 ; n25130_not
g36777 not n14060 ; n14060_not
g36778 not n12521 ; n12521_not
g36779 not n16112 ; n16112_not
g36780 not n15401 ; n15401_not
g36781 not n12611 ; n12611_not
g36782 not n26300 ; n26300_not
g36783 not n18011 ; n18011_not
g36784 not n11180 ; n11180_not
g36785 not n12440 ; n12440_not
g36786 not n10145 ; n10145_not
g36787 not n18110 ; n18110_not
g36788 not n16004 ; n16004_not
g36789 not n24023 ; n24023_not
g36790 not n23033 ; n23033_not
g36791 not n18002 ; n18002_not
g36792 not n20243 ; n20243_not
g36793 not n25112 ; n25112_not
g36794 not n21620 ; n21620_not
g36795 not n11153 ; n11153_not
g36796 not n20252 ; n20252_not
g36797 not n21215 ; n21215_not
g36798 not n20540 ; n20540_not
g36799 not n15311 ; n15311_not
g36800 not n23006 ; n23006_not
g36801 not n14213 ; n14213_not
g36802 not n12413 ; n12413_not
g36803 not n11162 ; n11162_not
g36804 not n25121 ; n25121_not
g36805 not n10127 ; n10127_not
g36806 not n16013 ; n16013_not
g36807 not n11144 ; n11144_not
g36808 not n23132 ; n23132_not
g36809 not n13340 ; n13340_not
g36810 not n17201 ; n17201_not
g36811 not n15131 ; n15131_not
g36812 not n10901 ; n10901_not
g36813 not n25103 ; n25103_not
g36814 not n10910 ; n10910_not
g36815 not n11171 ; n11171_not
g36816 not n20810 ; n20810_not
g36817 not n22241 ; n22241_not
g36818 not n22250 ; n22250_not
g36819 not n16103 ; n16103_not
g36820 not n16022 ; n16022_not
g36821 not n10064 ; n10064_not
g36822 not n14321 ; n14321_not
g36823 not n17012 ; n17012_not
g36824 not n24014 ; n24014_not
g36825 not n25301 ; n25301_not
g36826 not n17003 ; n17003_not
g36827 not n12008 ; n12008_not
g36828 not n22223 ; n22223_not
g36829 not n24032 ; n24032_not
g36830 not n11216 ; n11216_not
g36831 not n19010 ; n19010_not
g36832 not n13430 ; n13430_not
g36833 not n21008 ; n21008_not
g36834 not n10190 ; n10190_not
g36835 not n11072 ; n11072_not
g36836 not n10820 ; n10820_not
g36837 not n14051 ; n14051_not
g36838 not n15032 ; n15032_not
g36839 not n10244 ; n10244_not
g36840 not n20720 ; n20720_not
g36841 not n22340 ; n22340_not
g36842 not n22160 ; n22160_not
g36843 not n21206 ; n21206_not
g36844 not n16130 ; n16130_not
g36845 not n12053 ; n12053_not
g36846 not n21134 ; n21134_not
g36847 not n10046 ; n10046_not
g36848 not n10019 ; n10019_not
g36849 not n16031 ; n16031_not
g36850 not n10208 ; n10208_not
g36851 not n10217 ; n10217_not
g36852 not n20360 ; n20360_not
g36853 not n25004 ; n25004_not
g36854 not n22601 ; n22601_not
g36855 not n15113 ; n15113_not
g36856 not n10523 ; n10523_not
g36857 not n21170 ; n21170_not
g36858 not n10226 ; n10226_not
g36859 not n10235 ; n10235_not
g36860 not n11414 ; n11414_not
g36861 not n15023 ; n15023_not
g36862 not n27200 ; n27200_not
g36863 not n13304 ; n13304_not
g36864 not n14501 ; n14501_not
g36865 not n14033 ; n14033_not
g36866 not n13016 ; n13016_not
g36867 not n10802 ; n10802_not
g36868 not n14240 ; n14240_not
g36869 not n20180 ; n20180_not
g36870 not n11423 ; n11423_not
g36871 not n10262 ; n10262_not
g36872 not n14024 ; n14024_not
g36873 not n15014 ; n15014_not
g36874 not n14042 ; n14042_not
g36875 not n12062 ; n12062_not
g36876 not n21251 ; n21251_not
g36877 not n13421 ; n13421_not
g36878 not n12431 ; n12431_not
g36879 not n10253 ; n10253_not
g36880 not n11405 ; n11405_not
g36881 not n13601 ; n13601_not
g36882 not n10811 ; n10811_not
g36883 not n26003 ; n26003_not
g36884 not n14105 ; n14105_not
g36885 not n20351 ; n20351_not
g36886 not n21710 ; n21710_not
g36887 not n23150 ; n23150_not
g36888 not n27101 ; n27101_not
g36889 not n22322 ; n22322_not
g36890 not n11333 ; n11333_not
g36891 not n21350 ; n21350_not
g36892 not n11351 ; n11351_not
g36893 not n12503 ; n12503_not
g36894 not n20342 ; n20342_not
g36895 not n21143 ; n21143_not
g36896 not n24500 ; n24500_not
g36897 not n15050 ; n15050_not
g36898 not n14231 ; n14231_not
g36899 not n20054 ; n20054_not
g36900 not n13322 ; n13322_not
g36901 not n21341 ; n21341_not
g36902 not n22313 ; n22313_not
g36903 not n18020 ; n18020_not
g36904 not n21152 ; n21152_not
g36905 not n22331 ; n22331_not
g36906 not n11324 ; n11324_not
g36907 not n20270 ; n20270_not
g36908 not n22700 ; n22700_not
g36909 not n22304 ; n22304_not
g36910 not n11360 ; n11360_not
g36911 not n11108 ; n11108_not
g36912 not n12602 ; n12602_not
g36913 not n12108 ; n12108_not
g36914 not n23043 ; n23043_not
g36915 not n12063 ; n12063_not
g36916 not n15312 ; n15312_not
g36917 not n13305 ; n13305_not
g36918 not n12072 ; n12072_not
g36919 not n13332 ; n13332_not
g36920 not n23322 ; n23322_not
g36921 not n27102 ; n27102_not
g36922 not n25302 ; n25302_not
g36923 not n21027 ; n21027_not
g36924 not n12081 ; n12081_not
g36925 not n21621 ; n21621_not
g36926 not n20901 ; n20901_not
g36927 not n21531 ; n21531_not
g36928 not n13323 ; n13323_not
g36929 not n23160 ; n23160_not
g36930 not n12045 ; n12045_not
g36931 not n22710 ; n22710_not
g36932 not n13350 ; n13350_not
g36933 not n13341 ; n13341_not
g36934 not n12036 ; n12036_not
g36935 not n21630 ; n21630_not
g36936 not n23340 ; n23340_not
g36937 not n10515 ; n10515_not
g36938 not n21612 ; n21612_not
g36939 not n19020 ; n19020_not
g36940 not n21009 ; n21009_not
g36941 not n27003 ; n27003_not
g36942 not n10461 ; n10461_not
g36943 not n21018 ; n21018_not
g36944 not n20037 ; n20037_not
g36945 not n20055 ; n20055_not
g36946 not n12027 ; n12027_not
g36947 not n14223 ; n14223_not
g36948 not n20064 ; n20064_not
g36949 not n20046 ; n20046_not
g36950 not n10524 ; n10524_not
g36951 not n23313 ; n23313_not
g36952 not n13314 ; n13314_not
g36953 not n23331 ; n23331_not
g36954 not n14313 ; n14313_not
g36955 not n12018 ; n12018_not
g36956 not n12126 ; n12126_not
g36957 not n23304 ; n23304_not
g36958 not n12054 ; n12054_not
g36959 not n13260 ; n13260_not
g36960 not n12117 ; n12117_not
g36961 not n22413 ; n22413_not
g36962 not n15150 ; n15150_not
g36963 not n22701 ; n22701_not
g36964 not n21540 ; n21540_not
g36965 not n10533 ; n10533_not
g36966 not n10470 ; n10470_not
g36967 not n10506 ; n10506_not
g36968 not n13242 ; n13242_not
g36969 not n10173 ; n10173_not
g36970 not n21603 ; n21603_not
g36971 not n20910 ; n20910_not
g36972 not n12090 ; n12090_not
g36973 not n23412 ; n23412_not
g36974 not n12135 ; n12135_not
g36975 not n12009 ; n12009_not
g36976 not n13800 ; n13800_not
g36977 not n15204 ; n15204_not
g36978 not n10560 ; n10560_not
g36979 not n10542 ; n10542_not
g36980 not n21432 ; n21432_not
g36981 not n15600 ; n15600_not
g36982 not n21522 ; n21522_not
g36983 not n11712 ; n11712_not
g36984 not n27012 ; n27012_not
g36985 not n20073 ; n20073_not
g36986 not n21414 ; n21414_not
g36987 not n24600 ; n24600_not
g36988 not n12504 ; n12504_not
g36989 not n23151 ; n23151_not
g36990 not n21162 ; n21162_not
g36991 not n12513 ; n12513_not
g36992 not n15402 ; n15402_not
g36993 not n25032 ; n25032_not
g36994 not n12603 ; n12603_not
g36995 not n12522 ; n12522_not
g36996 not n21324 ; n21324_not
g36997 not n21171 ; n21171_not
g36998 not n10182 ; n10182_not
g36999 not n12531 ; n12531_not
g37000 not n15222 ; n15222_not
g37001 not n12900 ; n12900_not
g37002 not n23142 ; n23142_not
g37003 not n12540 ; n12540_not
g37004 not n25050 ; n25050_not
g37005 not n25041 ; n25041_not
g37006 not n21315 ; n21315_not
g37007 not n21180 ; n21180_not
g37008 not n22620 ; n22620_not
g37009 not n22800 ; n22800_not
g37010 not n21306 ; n21306_not
g37011 not n12252 ; n12252_not
g37012 not n12423 ; n12423_not
g37013 not n10254 ; n10254_not
g37014 not n12432 ; n12432_not
g37015 not n21117 ; n21117_not
g37016 not n15231 ; n15231_not
g37017 not n10245 ; n10245_not
g37018 not n25401 ; n25401_not
g37019 not n12450 ; n12450_not
g37020 not n10236 ; n10236_not
g37021 not n19101 ; n19101_not
g37022 not n10227 ; n10227_not
g37023 not n10218 ; n10218_not
g37024 not n21126 ; n21126_not
g37025 not n21360 ; n21360_not
g37026 not n10209 ; n10209_not
g37027 not n21135 ; n21135_not
g37028 not n15132 ; n15132_not
g37029 not n15042 ; n15042_not
g37030 not n15411 ; n15411_not
g37031 not n12207 ; n12207_not
g37032 not n25014 ; n25014_not
g37033 not n21144 ; n21144_not
g37034 not n15051 ; n15051_not
g37035 not n21342 ; n21342_not
g37036 not n21153 ; n21153_not
g37037 not n10191 ; n10191_not
g37038 not n25023 ; n25023_not
g37039 not n12630 ; n12630_not
g37040 not n10065 ; n10065_not
g37041 not n25131 ; n25131_not
g37042 not n10074 ; n10074_not
g37043 not n21225 ; n21225_not
g37044 not n25140 ; n25140_not
g37045 not n21270 ; n21270_not
g37046 not n21207 ; n21207_not
g37047 not n27300 ; n27300_not
g37048 not n17004 ; n17004_not
g37049 not n21252 ; n21252_not
g37050 not n15114 ; n15114_not
g37051 not n10092 ; n10092_not
g37052 not n23007 ; n23007_not
g37053 not n21234 ; n21234_not
g37054 not n17103 ; n17103_not
g37055 not n15123 ; n15123_not
g37056 not n25203 ; n25203_not
g37057 not n21243 ; n21243_not
g37058 not n25212 ; n25212_not
g37059 not n25221 ; n25221_not
g37060 not n12720 ; n12720_not
g37061 not n12621 ; n12621_not
g37062 not n12711 ; n12711_not
g37063 not n17130 ; n17130_not
g37064 not n17121 ; n17121_not
g37065 not n12702 ; n12702_not
g37066 not n17220 ; n17220_not
g37067 not n25320 ; n25320_not
g37068 not n10164 ; n10164_not
g37069 not n17211 ; n17211_not
g37070 not n17013 ; n17013_not
g37071 not n25104 ; n25104_not
g37072 not n25311 ; n25311_not
g37073 not n17202 ; n17202_not
g37074 not n23133 ; n23133_not
g37075 not n10155 ; n10155_not
g37076 not n17031 ; n17031_not
g37077 not n10056 ; n10056_not
g37078 not n25113 ; n25113_not
g37079 not n17040 ; n17040_not
g37080 not n15105 ; n15105_not
g37081 not n12612 ; n12612_not
g37082 not n12810 ; n12810_not
g37083 not n10128 ; n10128_not
g37084 not n12801 ; n12801_not
g37085 not n25122 ; n25122_not
g37086 not n21216 ; n21216_not
g37087 not n18210 ; n18210_not
g37088 not n12225 ; n12225_not
g37089 not n23232 ; n23232_not
g37090 not n27021 ; n27021_not
g37091 not n13143 ; n13143_not
g37092 not n21045 ; n21045_not
g37093 not n12243 ; n12243_not
g37094 not n13134 ; n13134_not
g37095 not n23214 ; n23214_not
g37096 not n12261 ; n12261_not
g37097 not n13125 ; n13125_not
g37098 not n20019 ; n20019_not
g37099 not n10371 ; n10371_not
g37100 not n13116 ; n13116_not
g37101 not n13008 ; n13008_not
g37102 not n23205 ; n23205_not
g37103 not n10362 ; n10362_not
g37104 not n21063 ; n21063_not
g37105 not n21072 ; n21072_not
g37106 not n13224 ; n13224_not
g37107 not n10380 ; n10380_not
g37108 not n10452 ; n10452_not
g37109 not n12153 ; n12153_not
g37110 not n20028 ; n20028_not
g37111 not n12162 ; n12162_not
g37112 not n13215 ; n13215_not
g37113 not n10443 ; n10443_not
g37114 not n13206 ; n13206_not
g37115 not n10416 ; n10416_not
g37116 not n12180 ; n12180_not
g37117 not n23250 ; n23250_not
g37118 not n15501 ; n15501_not
g37119 not n24510 ; n24510_not
g37120 not n10434 ; n10434_not
g37121 not n21504 ; n21504_not
g37122 not n10425 ; n10425_not
g37123 not n13170 ; n13170_not
g37124 not n17400 ; n17400_not
g37125 not n15321 ; n15321_not
g37126 not n10407 ; n10407_not
g37127 not n13161 ; n13161_not
g37128 not n15141 ; n15141_not
g37129 not n23241 ; n23241_not
g37130 not n12216 ; n12216_not
g37131 not n13053 ; n13053_not
g37132 not n12351 ; n12351_not
g37133 not n20550 ; n20550_not
g37134 not n21423 ; n21423_not
g37135 not n23106 ; n23106_not
g37136 not n17310 ; n17310_not
g37137 not n25410 ; n25410_not
g37138 not n15006 ; n15006_not
g37139 not n10038 ; n10038_not
g37140 not n13026 ; n13026_not
g37141 not n17301 ; n17301_not
g37142 not n20820 ; n20820_not
g37143 not n10281 ; n10281_not
g37144 not n15420 ; n15420_not
g37145 not n12405 ; n12405_not
g37146 not n15015 ; n15015_not
g37147 not n10272 ; n10272_not
g37148 not n12315 ; n12315_not
g37149 not n13017 ; n13017_not
g37150 not n10263 ; n10263_not
g37151 not n21108 ; n21108_not
g37152 not n15303 ; n15303_not
g37153 not n15024 ; n15024_not
g37154 not n13107 ; n13107_not
g37155 not n10344 ; n10344_not
g37156 not n22602 ; n22602_not
g37157 not n12306 ; n12306_not
g37158 not n10326 ; n10326_not
g37159 not n10317 ; n10317_not
g37160 not n12324 ; n12324_not
g37161 not n15213 ; n15213_not
g37162 not n10308 ; n10308_not
g37163 not n21081 ; n21081_not
g37164 not n21450 ; n21450_not
g37165 not n21441 ; n21441_not
g37166 not n12342 ; n12342_not
g37167 not n13080 ; n13080_not
g37168 not n21090 ; n21090_not
g37169 not n10029 ; n10029_not
g37170 not n13044 ; n13044_not
g37171 not n13071 ; n13071_not
g37172 not n12360 ; n12360_not
g37173 not n13062 ; n13062_not
g37174 not n19110 ; n19110_not
g37175 not n27030 ; n27030_not
g37176 not n11622 ; n11622_not
g37177 not n14421 ; n14421_not
g37178 not n20523 ; n20523_not
g37179 not n22314 ; n22314_not
g37180 not n20118 ; n20118_not
g37181 not n22170 ; n22170_not
g37182 not n11631 ; n11631_not
g37183 not n23052 ; n23052_not
g37184 not n22107 ; n22107_not
g37185 not n23124 ; n23124_not
g37186 not n11280 ; n11280_not
g37187 not n20109 ; n20109_not
g37188 not n14133 ; n14133_not
g37189 not n24231 ; n24231_not
g37190 not n11640 ; n11640_not
g37191 not n20244 ; n20244_not
g37192 not n26121 ; n26121_not
g37193 not n24240 ; n24240_not
g37194 not n20532 ; n20532_not
g37195 not n11271 ; n11271_not
g37196 not n16122 ; n16122_not
g37197 not n22125 ; n22125_not
g37198 not n24042 ; n24042_not
g37199 not n20145 ; n20145_not
g37200 not n20226 ; n20226_not
g37201 not n14430 ; n14430_not
g37202 not n10713 ; n10713_not
g37203 not n22422 ; n22422_not
g37204 not n24204 ; n24204_not
g37205 not n20505 ; n20505_not
g37206 not n22440 ; n22440_not
g37207 not n14115 ; n14115_not
g37208 not n22116 ; n22116_not
g37209 not n26130 ; n26130_not
g37210 not n10704 ; n10704_not
g37211 not n14610 ; n14610_not
g37212 not n24015 ; n24015_not
g37213 not n24213 ; n24213_not
g37214 not n20136 ; n20136_not
g37215 not n11604 ; n11604_not
g37216 not n20127 ; n20127_not
g37217 not n20514 ; n20514_not
g37218 not n11613 ; n11613_not
g37219 not n24222 ; n24222_not
g37220 not n24312 ; n24312_not
g37221 not n14160 ; n14160_not
g37222 not n22260 ; n22260_not
g37223 not n11703 ; n11703_not
g37224 not n22062 ; n22062_not
g37225 not n11235 ; n11235_not
g37226 not n24321 ; n24321_not
g37227 not n11109 ; n11109_not
g37228 not n20235 ; n20235_not
g37229 not n11307 ; n11307_not
g37230 not n22512 ; n22512_not
g37231 not n10650 ; n10650_not
g37232 not n22071 ; n22071_not
g37233 not n10902 ; n10902_not
g37234 not n11721 ; n11721_not
g37235 not n22053 ; n22053_not
g37236 not n24330 ; n24330_not
g37237 not n11226 ; n11226_not
g37238 not n11325 ; n11325_not
g37239 not n10911 ; n10911_not
g37240 not n15330 ; n15330_not
g37241 not n23520 ; n23520_not
g37242 not n22242 ; n22242_not
g37243 not n16302 ; n16302_not
g37244 not n20325 ; n20325_not
g37245 not n14142 ; n14142_not
g37246 not n22503 ; n22503_not
g37247 not n22080 ; n22080_not
g37248 not n11262 ; n11262_not
g37249 not n16311 ; n16311_not
g37250 not n16113 ; n16113_not
g37251 not n16320 ; n16320_not
g37252 not n14151 ; n14151_not
g37253 not n26112 ; n26112_not
g37254 not n14412 ; n14412_not
g37255 not n24303 ; n24303_not
g37256 not n26103 ; n26103_not
g37257 not n10353 ; n10353_not
g37258 not n14403 ; n14403_not
g37259 not n11244 ; n11244_not
g37260 not n23016 ; n23016_not
g37261 not n14025 ; n14025_not
g37262 not n11406 ; n11406_not
g37263 not n20361 ; n20361_not
g37264 not n11370 ; n11370_not
g37265 not n14502 ; n14502_not
g37266 not n11433 ; n11433_not
g37267 not n14016 ; n14016_not
g37268 not n16131 ; n16131_not
g37269 not n14205 ; n14205_not
g37270 not n14511 ; n14511_not
g37271 not n22332 ; n22332_not
g37272 not n10821 ; n10821_not
g37273 not n11451 ; n11451_not
g37274 not n23700 ; n23700_not
g37275 not n20406 ; n20406_not
g37276 not n24060 ; n24060_not
g37277 not n11361 ; n11361_not
g37278 not n26202 ; n26202_not
g37279 not n14520 ; n14520_not
g37280 not n20172 ; n20172_not
g37281 not n18201 ; n18201_not
g37282 not n19011 ; n19011_not
g37283 not n27201 ; n27201_not
g37284 not n22323 ; n22323_not
g37285 not n10830 ; n10830_not
g37286 not n20352 ; n20352_not
g37287 not n14061 ; n14061_not
g37288 not n14052 ; n14052_not
g37289 not n22044 ; n22044_not
g37290 not n14070 ; n14070_not
g37291 not n22341 ; n22341_not
g37292 not n26211 ; n26211_not
g37293 not n14043 ; n14043_not
g37294 not n16140 ; n16140_not
g37295 not n13611 ; n13611_not
g37296 not n10812 ; n10812_not
g37297 not n20370 ; n20370_not
g37298 not n14034 ; n14034_not
g37299 not n20181 ; n20181_not
g37300 not n11415 ; n11415_not
g37301 not n10803 ; n10803_not
g37302 not n11523 ; n11523_not
g37303 not n24123 ; n24123_not
g37304 not n27120 ; n27120_not
g37305 not n24132 ; n24132_not
g37306 not n22305 ; n22305_not
g37307 not n14106 ; n14106_not
g37308 not n11532 ; n11532_not
g37309 not n20451 ; n20451_not
g37310 not n10731 ; n10731_not
g37311 not n16212 ; n16212_not
g37312 not n11541 ; n11541_not
g37313 not n20208 ; n20208_not
g37314 not n24141 ; n24141_not
g37315 not n22431 ; n22431_not
g37316 not n20460 ; n20460_not
g37317 not n11316 ; n11316_not
g37318 not n16221 ; n16221_not
g37319 not n11550 ; n11550_not
g37320 not n20217 ; n20217_not
g37321 not n22134 ; n22134_not
g37322 not n23601 ; n23601_not
g37323 not n16230 ; n16230_not
g37324 not n14601 ; n14601_not
g37325 not n13521 ; n13521_not
g37326 not n22143 ; n22143_not
g37327 not n22404 ; n22404_not
g37328 not n22251 ; n22251_not
g37329 not n20163 ; n20163_not
g37330 not n11352 ; n11352_not
g37331 not n20424 ; n20424_not
g37332 not n24105 ; n24105_not
g37333 not n20433 ; n20433_not
g37334 not n23502 ; n23502_not
g37335 not n24051 ; n24051_not
g37336 not n24114 ; n24114_not
g37337 not n26220 ; n26220_not
g37338 not n20190 ; n20190_not
g37339 not n11505 ; n11505_not
g37340 not n11343 ; n11343_not
g37341 not n20343 ; n20343_not
g37342 not n23610 ; n23610_not
g37343 not n20442 ; n20442_not
g37344 not n20154 ; n20154_not
g37345 not n20262 ; n20262_not
g37346 not n18030 ; n18030_not
g37347 not n16500 ; n16500_not
g37348 not n20721 ; n20721_not
g37349 not n11118 ; n11118_not
g37350 not n19002 ; n19002_not
g37351 not n26310 ; n26310_not
g37352 not n20730 ; n20730_not
g37353 not n20271 ; n20271_not
g37354 not n21810 ; n21810_not
g37355 not n14232 ; n14232_not
g37356 not n24501 ; n24501_not
g37357 not n26301 ; n26301_not
g37358 not n16032 ; n16032_not
g37359 not n20640 ; n20640_not
g37360 not n13530 ; n13530_not
g37361 not n21801 ; n21801_not
g37362 not n14304 ; n14304_not
g37363 not n24411 ; n24411_not
g37364 not n26013 ; n26013_not
g37365 not n16023 ; n16023_not
g37366 not n21900 ; n21900_not
g37367 not n24420 ; n24420_not
g37368 not n14214 ; n14214_not
g37369 not n23421 ; n23421_not
g37370 not n11154 ; n11154_not
g37371 not n20703 ; n20703_not
g37372 not n18021 ; n18021_not
g37373 not n13620 ; n13620_not
g37374 not n14331 ; n14331_not
g37375 not n11145 ; n11145_not
g37376 not n18102 ; n18102_not
g37377 not n26004 ; n26004_not
g37378 not n20712 ; n20712_not
g37379 not n11136 ; n11136_not
g37380 not n13602 ; n13602_not
g37381 not n20091 ; n20091_not
g37382 not n16203 ; n16203_not
g37383 not n20253 ; n20253_not
g37384 not n16050 ; n16050_not
g37385 not n21720 ; n21720_not
g37386 not n11055 ; n11055_not
g37387 not n21711 ; n21711_not
g37388 not n23430 ; n23430_not
g37389 not n13431 ; n13431_not
g37390 not n23115 ; n23115_not
g37391 not n19200 ; n19200_not
g37392 not n11046 ; n11046_not
g37393 not n11019 ; n11019_not
g37394 not n22215 ; n22215_not
g37395 not n13422 ; n13422_not
g37396 not n20082 ; n20082_not
g37397 not n21702 ; n21702_not
g37398 not n11037 ; n11037_not
g37399 not n23034 ; n23034_not
g37400 not n13413 ; n13413_not
g37401 not n11028 ; n11028_not
g37402 not n27111 ; n27111_not
g37403 not n20802 ; n20802_not
g37404 not n23061 ; n23061_not
g37405 not n14241 ; n14241_not
g37406 not n11901 ; n11901_not
g37407 not n11091 ; n11091_not
g37408 not n20307 ; n20307_not
g37409 not n20280 ; n20280_not
g37410 not n13503 ; n13503_not
g37411 not n11082 ; n11082_not
g37412 not n22611 ; n22611_not
g37413 not n22206 ; n22206_not
g37414 not n11073 ; n11073_not
g37415 not n11910 ; n11910_not
g37416 not n20811 ; n20811_not
g37417 not n24006 ; n24006_not
g37418 not n23070 ; n23070_not
g37419 not n14250 ; n14250_not
g37420 not n16041 ; n16041_not
g37421 not n20541 ; n20541_not
g37422 not n18111 ; n18111_not
g37423 not n11181 ; n11181_not
g37424 not n23511 ; n23511_not
g37425 not n26040 ; n26040_not
g37426 not n18012 ; n18012_not
g37427 not n22017 ; n22017_not
g37428 not n22224 ; n22224_not
g37429 not n13710 ; n13710_not
g37430 not n26031 ; n26031_not
g37431 not n24402 ; n24402_not
g37432 not n11172 ; n11172_not
g37433 not n23025 ; n23025_not
g37434 not n16014 ; n16014_not
g37435 not n22008 ; n22008_not
g37436 not n11208 ; n11208_not
g37437 not n26022 ; n26022_not
g37438 not n10740 ; n10740_not
g37439 not n22035 ; n22035_not
g37440 not n10623 ; n10623_not
g37441 not n10920 ; n10920_not
g37442 not n16401 ; n16401_not
g37443 not n18120 ; n18120_not
g37444 not n18003 ; n18003_not
g37445 not n11190 ; n11190_not
g37446 not n10632 ; n10632_not
g37447 not n20631 ; n20631_not
g37448 not n20622 ; n20622_not
g37449 not n13701 ; n13701_not
g37450 not n16410 ; n16410_not
g37451 not n24024 ; n24024_not
g37452 not n16005 ; n16005_not
g37453 not n20316 ; n20316_not
g37454 not n20613 ; n20613_not
g37455 not n10614 ; n10614_not
g37456 not n11217 ; n11217_not
g37457 not n11442 ; n11442_not
g37458 not n10641 ; n10641_not
g37459 not n10605 ; n10605_not
g37460 not n11811 ; n11811_not
g37461 not n22521 ; n22521_not
g37462 not n11730 ; n11730_not
g37463 not n24033 ; n24033_not
g37464 not n11802 ; n11802_not
g37465 not n17122 ; n17122_not
g37466 not n22225 ; n22225_not
g37467 not n14251 ; n14251_not
g37468 not n22171 ; n22171_not
g37469 not n17023 ; n17023_not
g37470 not n14161 ; n14161_not
g37471 not n14071 ; n14071_not
g37472 not n22324 ; n22324_not
g37473 not n14170 ; n14170_not
g37474 not n24070 ; n24070_not
g37475 not n22243 ; n22243_not
g37476 not n22234 ; n22234_not
g37477 not n15124 ; n15124_not
g37478 not n25015 ; n25015_not
g37479 not n14080 ; n14080_not
g37480 not n21181 ; n21181_not
g37481 not n17104 ; n17104_not
g37482 not n16033 ; n16033_not
g37483 not n17014 ; n17014_not
g37484 not n13207 ; n13207_not
g37485 not n23134 ; n23134_not
g37486 not n14062 ; n14062_not
g37487 not n12712 ; n12712_not
g37488 not n12703 ; n12703_not
g37489 not n17032 ; n17032_not
g37490 not n16105 ; n16105_not
g37491 not n12721 ; n12721_not
g37492 not n16051 ; n16051_not
g37493 not n16141 ; n16141_not
g37494 not n25213 ; n25213_not
g37495 not n21361 ; n21361_not
g37496 not n22180 ; n22180_not
g37497 not n16150 ; n16150_not
g37498 not n22333 ; n22333_not
g37499 not n16132 ; n16132_not
g37500 not n15412 ; n15412_not
g37501 not n21370 ; n21370_not
g37502 not n22207 ; n22207_not
g37503 not n12730 ; n12730_not
g37504 not n14260 ; n14260_not
g37505 not n25204 ; n25204_not
g37506 not n23116 ; n23116_not
g37507 not n16042 ; n16042_not
g37508 not n25105 ; n25105_not
g37509 not n24061 ; n24061_not
g37510 not n12406 ; n12406_not
g37511 not n25033 ; n25033_not
g37512 not n14107 ; n14107_not
g37513 not n14116 ; n14116_not
g37514 not n21316 ; n21316_not
g37515 not n14134 ; n14134_not
g37516 not n17050 ; n17050_not
g37517 not n25051 ; n25051_not
g37518 not n15106 ; n15106_not
g37519 not n16024 ; n16024_not
g37520 not n12811 ; n12811_not
g37521 not n23053 ; n23053_not
g37522 not n14314 ; n14314_not
g37523 not n23062 ; n23062_not
g37524 not n25132 ; n25132_not
g37525 not n14440 ; n14440_not
g37526 not n14224 ; n14224_not
g37527 not n14143 ; n14143_not
g37528 not n23143 ; n23143_not
g37529 not n16015 ; n16015_not
g37530 not n16123 ; n16123_not
g37531 not n22900 ; n22900_not
g37532 not n12802 ; n12802_not
g37533 not n16006 ; n16006_not
g37534 not n17041 ; n17041_not
g37535 not n14422 ; n14422_not
g37536 not n24043 ; n24043_not
g37537 not n14215 ; n14215_not
g37538 not n14125 ; n14125_not
g37539 not n24016 ; n24016_not
g37540 not n25123 ; n25123_not
g37541 not n14332 ; n14332_not
g37542 not n15331 ; n15331_not
g37543 not n21325 ; n21325_not
g37544 not n14431 ; n14431_not
g37545 not n25042 ; n25042_not
g37546 not n23800 ; n23800_not
g37547 not n21253 ; n21253_not
g37548 not n23620 ; n23620_not
g37549 not n15052 ; n15052_not
g37550 not n25024 ; n25024_not
g37551 not n14233 ; n14233_not
g37552 not n14404 ; n14404_not
g37553 not n16060 ; n16060_not
g37554 not n24025 ; n24025_not
g37555 not n14242 ; n14242_not
g37556 not n16114 ; n16114_not
g37557 not n22315 ; n22315_not
g37558 not n15223 ; n15223_not
g37559 not n22153 ; n22153_not
g37560 not n25114 ; n25114_not
g37561 not n22261 ; n22261_not
g37562 not n21343 ; n21343_not
g37563 not n24052 ; n24052_not
g37564 not n24007 ; n24007_not
g37565 not n14350 ; n14350_not
g37566 not n15061 ; n15061_not
g37567 not n25060 ; n25060_not
g37568 not n21307 ; n21307_not
g37569 not n15403 ; n15403_not
g37570 not n21334 ; n21334_not
g37571 not n25141 ; n25141_not
g37572 not n21271 ; n21271_not
g37573 not n23035 ; n23035_not
g37574 not n15322 ; n15322_not
g37575 not n25150 ; n25150_not
g37576 not n12820 ; n12820_not
g37577 not n23152 ; n23152_not
g37578 not n14413 ; n14413_not
g37579 not n22306 ; n22306_not
g37580 not n21262 ; n21262_not
g37581 not n13630 ; n13630_not
g37582 not n21460 ; n21460_not
g37583 not n21550 ; n21550_not
g37584 not n21541 ; n21541_not
g37585 not n15700 ; n15700_not
g37586 not n23323 ; n23323_not
g37587 not n23125 ; n23125_not
g37588 not n23080 ; n23080_not
g37589 not n22009 ; n22009_not
g37590 not n22540 ; n22540_not
g37591 not n14710 ; n14710_not
g37592 not n22531 ; n22531_not
g37593 not n24403 ; n24403_not
g37594 not n22522 ; n22522_not
g37595 not n23161 ; n23161_not
g37596 not n23314 ; n23314_not
g37597 not n23341 ; n23341_not
g37598 not n13306 ; n13306_not
g37599 not n24430 ; n24430_not
g37600 not n16501 ; n16501_not
g37601 not n21901 ; n21901_not
g37602 not n23422 ; n23422_not
g37603 not n22702 ; n22702_not
g37604 not n13612 ; n13612_not
g37605 not n22711 ; n22711_not
g37606 not n13621 ; n13621_not
g37607 not n24421 ; n24421_not
g37608 not n23332 ; n23332_not
g37609 not n15205 ; n15205_not
g37610 not n21604 ; n21604_not
g37611 not n13234 ; n13234_not
g37612 not n23512 ; n23512_not
g37613 not n13225 ; n13225_not
g37614 not n22036 ; n22036_not
g37615 not n24340 ; n24340_not
g37616 not n15520 ; n15520_not
g37617 not n13720 ; n13720_not
g37618 not n15151 ; n15151_not
g37619 not n23260 ; n23260_not
g37620 not n24106 ; n24106_not
g37621 not n22801 ; n22801_not
g37622 not n13216 ; n13216_not
g37623 not n15502 ; n15502_not
g37624 not n23521 ; n23521_not
g37625 not n16420 ; n16420_not
g37626 not n22018 ; n22018_not
g37627 not n23026 ; n23026_not
g37628 not n21523 ; n21523_not
g37629 not n16411 ; n16411_not
g37630 not n24232 ; n24232_not
g37631 not n15340 ; n15340_not
g37632 not n13423 ; n13423_not
g37633 not n13243 ; n13243_not
g37634 not n16402 ; n16402_not
g37635 not n23305 ; n23305_not
g37636 not n22027 ; n22027_not
g37637 not n13702 ; n13702_not
g37638 not n27301 ; n27301_not
g37639 not n23044 ; n23044_not
g37640 not n13351 ; n13351_not
g37641 not n21622 ; n21622_not
g37642 not n23224 ; n23224_not
g37643 not n13450 ; n13450_not
g37644 not n21721 ; n21721_not
g37645 not n13342 ; n13342_not
g37646 not n22630 ; n22630_not
g37647 not n13333 ; n13333_not
g37648 not n15241 ; n15241_not
g37649 not n15250 ; n15250_not
g37650 not n23431 ; n23431_not
g37651 not n23071 ; n23071_not
g37652 not n23404 ; n23404_not
g37653 not n16312 ; n16312_not
g37654 not n21730 ; n21730_not
g37655 not n13405 ; n13405_not
g37656 not n15313 ; n15313_not
g37657 not n23413 ; n23413_not
g37658 not n22621 ; n22621_not
g37659 not n13414 ; n13414_not
g37660 not n24601 ; n24601_not
g37661 not n21640 ; n21640_not
g37662 not n21703 ; n21703_not
g37663 not n21631 ; n21631_not
g37664 not n24610 ; n24610_not
g37665 not n13432 ; n13432_not
g37666 not n13360 ; n13360_not
g37667 not n22603 ; n22603_not
g37668 not n21613 ; n21613_not
g37669 not n15304 ; n15304_not
g37670 not n21802 ; n21802_not
g37671 not n13531 ; n13531_not
g37672 not n24502 ; n24502_not
g37673 not n13540 ; n13540_not
g37674 not n13324 ; n13324_not
g37675 not n21811 ; n21811_not
g37676 not n21820 ; n21820_not
g37677 not n21712 ; n21712_not
g37678 not n13315 ; n13315_not
g37679 not n16510 ; n16510_not
g37680 not n24511 ; n24511_not
g37681 not n24520 ; n24520_not
g37682 not n16600 ; n16600_not
g37683 not n22612 ; n22612_not
g37684 not n14800 ; n14800_not
g37685 not n15610 ; n15610_not
g37686 not n13504 ; n13504_not
g37687 not n24331 ; n24331_not
g37688 not n23440 ; n23440_not
g37689 not n15214 ; n15214_not
g37690 not n13522 ; n13522_not
g37691 not n15601 ; n15601_not
g37692 not n23350 ; n23350_not
g37693 not n13072 ; n13072_not
g37694 not n23611 ; n23611_not
g37695 not n22423 ; n22423_not
g37696 not n13063 ; n13063_not
g37697 not n21424 ; n21424_not
g37698 not n24115 ; n24115_not
g37699 not n13054 ; n13054_not
g37700 not n22414 ; n22414_not
g37701 not n13045 ; n13045_not
g37702 not n22405 ; n22405_not
g37703 not n22144 ; n22144_not
g37704 not n22135 ; n22135_not
g37705 not n15430 ; n15430_not
g37706 not n22126 ; n22126_not
g37707 not n24160 ; n24160_not
g37708 not n16231 ; n16231_not
g37709 not n24151 ; n24151_not
g37710 not n24142 ; n24142_not
g37711 not n23602 ; n23602_not
g37712 not n16213 ; n16213_not
g37713 not n13090 ; n13090_not
g37714 not n21442 ; n21442_not
g37715 not n16204 ; n16204_not
g37716 not n21433 ; n21433_not
g37717 not n24133 ; n24133_not
g37718 not n13081 ; n13081_not
g37719 not n24124 ; n24124_not
g37720 not n15133 ; n15133_not
g37721 not n22342 ; n22342_not
g37722 not n14035 ; n14035_not
g37723 not n13009 ; n13009_not
g37724 not n21154 ; n21154_not
g37725 not n15025 ; n15025_not
g37726 not n14206 ; n14206_not
g37727 not n15232 ; n15232_not
g37728 not n21406 ; n21406_not
g37729 not n14044 ; n14044_not
g37730 not n22162 ; n22162_not
g37731 not n14053 ; n14053_not
g37732 not n22252 ; n22252_not
g37733 not n15007 ; n15007_not
g37734 not n13027 ; n13027_not
g37735 not n14530 ; n14530_not
g37736 not n22360 ; n22360_not
g37737 not n23701 ; n23701_not
g37738 not n15421 ; n15421_not
g37739 not n14521 ; n14521_not
g37740 not n22351 ; n22351_not
g37741 not n14017 ; n14017_not
g37742 not n13018 ; n13018_not
g37743 not n14503 ; n14503_not
g37744 not n15016 ; n15016_not
g37745 not n23710 ; n23710_not
g37746 not n23242 ; n23242_not
g37747 not n21235 ; n21235_not
g37748 not n24304 ; n24304_not
g37749 not n22504 ; n22504_not
g37750 not n13162 ; n13162_not
g37751 not n22072 ; n22072_not
g37752 not n16330 ; n16330_not
g37753 not n16321 ; n16321_not
g37754 not n13153 ; n13153_not
g37755 not n22081 ; n22081_not
g37756 not n22054 ; n22054_not
g37757 not n22045 ; n22045_not
g37758 not n24322 ; n24322_not
g37759 not n24700 ; n24700_not
g37760 not n23530 ; n23530_not
g37761 not n22063 ; n22063_not
g37762 not n21505 ; n21505_not
g37763 not n13180 ; n13180_not
g37764 not n22513 ; n22513_not
g37765 not n23251 ; n23251_not
g37766 not n24313 ; n24313_not
g37767 not n21226 ; n21226_not
g37768 not n27310 ; n27310_not
g37769 not n15160 ; n15160_not
g37770 not n22108 ; n22108_not
g37771 not n24223 ; n24223_not
g37772 not n23017 ; n23017_not
g37773 not n15043 ; n15043_not
g37774 not n24214 ; n24214_not
g37775 not n22450 ; n22450_not
g37776 not n14620 ; n14620_not
g37777 not n13108 ; n13108_not
g37778 not n22441 ; n22441_not
g37779 not n14602 ; n14602_not
g37780 not n13900 ; n13900_not
g37781 not n24250 ; n24250_not
g37782 not n13801 ; n13801_not
g37783 not n16303 ; n16303_not
g37784 not n23233 ; n23233_not
g37785 not n13135 ; n13135_not
g37786 not n13144 ; n13144_not
g37787 not n13810 ; n13810_not
g37788 not n24241 ; n24241_not
g37789 not n22090 ; n22090_not
g37790 not n23206 ; n23206_not
g37791 not n23215 ; n23215_not
g37792 not n13117 ; n13117_not
g37793 not n13126 ; n13126_not
g37794 not n12280 ; n12280_not
g37795 not n10219 ; n10219_not
g37796 not n10228 ; n10228_not
g37797 not n10237 ; n10237_not
g37798 not n12262 ; n12262_not
g37799 not n11560 ; n11560_not
g37800 not n20173 ; n20173_not
g37801 not n20164 ; n20164_not
g37802 not n21046 ; n21046_not
g37803 not n12244 ; n12244_not
g37804 not n10507 ; n10507_not
g37805 not n10255 ; n10255_not
g37806 not n12235 ; n12235_not
g37807 not n26131 ; n26131_not
g37808 not n18220 ; n18220_not
g37809 not n20317 ; n20317_not
g37810 not n20452 ; n20452_not
g37811 not n12343 ; n12343_not
g37812 not n21082 ; n21082_not
g37813 not n10066 ; n10066_not
g37814 not n11542 ; n11542_not
g37815 not n10183 ; n10183_not
g37816 not n20461 ; n20461_not
g37817 not n12334 ; n12334_not
g37818 not n11551 ; n11551_not
g37819 not n12325 ; n12325_not
g37820 not n12307 ; n12307_not
g37821 not n20470 ; n20470_not
g37822 not n10192 ; n10192_not
g37823 not n19210 ; n19210_not
g37824 not n21064 ; n21064_not
g37825 not n26041 ; n26041_not
g37826 not n12190 ; n12190_not
g37827 not n11632 ; n11632_not
g37828 not n11641 ; n11641_not
g37829 not n26122 ; n26122_not
g37830 not n11650 ; n11650_not
g37831 not n27031 ; n27031_not
g37832 not n21037 ; n21037_not
g37833 not n17410 ; n17410_not
g37834 not n10318 ; n10318_not
g37835 not n12181 ; n12181_not
g37836 not n20155 ; n20155_not
g37837 not n17401 ; n17401_not
g37838 not n10732 ; n10732_not
g37839 not n12145 ; n12145_not
g37840 not n10750 ; n10750_not
g37841 not n12226 ; n12226_not
g37842 not n20506 ; n20506_not
g37843 not n10264 ; n10264_not
g37844 not n20227 ; n20227_not
g37845 not n20515 ; n20515_not
g37846 not n12208 ; n12208_not
g37847 not n10273 ; n10273_not
g37848 not n11614 ; n11614_not
g37849 not n20524 ; n20524_not
g37850 not n11623 ; n11623_not
g37851 not n10282 ; n10282_not
g37852 not n20191 ; n20191_not
g37853 not n10831 ; n10831_not
g37854 not n12451 ; n12451_not
g37855 not n25402 ; n25402_not
g37856 not n11425 ; n11425_not
g37857 not n12442 ; n12442_not
g37858 not n10822 ; n10822_not
g37859 not n11434 ; n11434_not
g37860 not n21118 ; n21118_not
g37861 not n10093 ; n10093_not
g37862 not n20074 ; n20074_not
g37863 not n11452 ; n11452_not
g37864 not n26203 ; n26203_not
g37865 not n20407 ; n20407_not
g37866 not n11461 ; n11461_not
g37867 not n12433 ; n12433_not
g37868 not n11083 ; n11083_not
g37869 not n26500 ; n26500_not
g37870 not n20380 ; n20380_not
g37871 not n21136 ; n21136_not
g37872 not n12037 ; n12037_not
g37873 not n12460 ; n12460_not
g37874 not n10039 ; n10039_not
g37875 not n26212 ; n26212_not
g37876 not n21127 ; n21127_not
g37877 not n10840 ; n10840_not
g37878 not n10057 ; n10057_not
g37879 not n12019 ; n12019_not
g37880 not n11407 ; n11407_not
g37881 not n11416 ; n11416_not
g37882 not n10075 ; n10075_not
g37883 not n11371 ; n11371_not
g37884 not n11362 ; n11362_not
g37885 not n10156 ; n10156_not
g37886 not n11290 ; n11290_not
g37887 not n25420 ; n25420_not
g37888 not n10165 ; n10165_not
g37889 not n20425 ; n20425_not
g37890 not n12370 ; n12370_not
g37891 not n20182 ; n20182_not
g37892 not n11506 ; n11506_not
g37893 not n12361 ; n12361_not
g37894 not n10174 ; n10174_not
g37895 not n10804 ; n10804_not
g37896 not n20443 ; n20443_not
g37897 not n18211 ; n18211_not
g37898 not n11524 ; n11524_not
g37899 not n12352 ; n12352_not
g37900 not n12424 ; n12424_not
g37901 not n18202 ; n18202_not
g37902 not n12415 ; n12415_not
g37903 not n21109 ; n21109_not
g37904 not n11470 ; n11470_not
g37905 not n12316 ; n12316_not
g37906 not n27040 ; n27040_not
g37907 not n10129 ; n10129_not
g37908 not n17302 ; n17302_not
g37909 not n10138 ; n10138_not
g37910 not n20416 ; n20416_not
g37911 not n10147 ; n10147_not
g37912 not n25411 ; n25411_not
g37913 not n17311 ; n17311_not
g37914 not n26023 ; n26023_not
g37915 not n11443 ; n11443_not
g37916 not n11803 ; n11803_not
g37917 not n11812 ; n11812_not
g37918 not n20911 ; n20911_not
g37919 not n20038 ; n20038_not
g37920 not n26014 ; n26014_not
g37921 not n20902 ; n20902_not
g37922 not n10615 ; n10615_not
g37923 not n10471 ; n10471_not
g37924 not n27004 ; n27004_not
g37925 not n20614 ; n20614_not
g37926 not n10480 ; n10480_not
g37927 not n10444 ; n10444_not
g37928 not n20623 ; n20623_not
g37929 not n10642 ; n10642_not
g37930 not n20704 ; n20704_not
g37931 not n10651 ; n10651_not
g37932 not n20920 ; n20920_not
g37933 not n20029 ; n20029_not
g37934 not n26050 ; n26050_not
g37935 not n25600 ; n25600_not
g37936 not n10453 ; n10453_not
g37937 not n10633 ; n10633_not
g37938 not n10624 ; n10624_not
g37939 not n20641 ; n20641_not
g37940 not n26032 ; n26032_not
g37941 not n20650 ; n20650_not
g37942 not n18310 ; n18310_not
g37943 not n10525 ; n10525_not
g37944 not n10534 ; n10534_not
g37945 not n20083 ; n20083_not
g37946 not n20740 ; n20740_not
g37947 not n10543 ; n10543_not
g37948 not n11920 ; n11920_not
g37949 not n20812 ; n20812_not
g37950 not n10561 ; n10561_not
g37951 not n11911 ; n11911_not
g37952 not n10552 ; n10552_not
g37953 not n20803 ; n20803_not
g37954 not n11902 ; n11902_not
g37955 not n20065 ; n20065_not
g37956 not n11830 ; n11830_not
g37957 not n10606 ; n10606_not
g37958 not n17320 ; n17320_not
g37959 not n26005 ; n26005_not
g37960 not n20047 ; n20047_not
g37961 not n20830 ; n20830_not
g37962 not n20713 ; n20713_not
g37963 not n10516 ; n10516_not
g37964 not n20092 ; n20092_not
g37965 not n20821 ; n20821_not
g37966 not n20722 ; n20722_not
g37967 not n10705 ; n10705_not
g37968 not n10363 ; n10363_not
g37969 not n12127 ; n12127_not
g37970 not n26104 ; n26104_not
g37971 not n20542 ; n20542_not
g37972 not n12118 ; n12118_not
g37973 not n20551 ; n20551_not
g37974 not n20137 ; n20137_not
g37975 not n12109 ; n12109_not
g37976 not n20560 ; n20560_not
g37977 not n11704 ; n11704_not
g37978 not n10381 ; n10381_not
g37979 not n20533 ; n20533_not
g37980 not n25510 ; n25510_not
g37981 not n10327 ; n10327_not
g37982 not n12163 ; n12163_not
g37983 not n12154 ; n12154_not
g37984 not n26113 ; n26113_not
g37985 not n21028 ; n21028_not
g37986 not n10336 ; n10336_not
g37987 not n10723 ; n10723_not
g37988 not n10345 ; n10345_not
g37989 not n12136 ; n12136_not
g37990 not n11731 ; n11731_not
g37991 not n12073 ; n12073_not
g37992 not n18400 ; n18400_not
g37993 not n11740 ; n11740_not
g37994 not n10660 ; n10660_not
g37995 not n12055 ; n12055_not
g37996 not n18004 ; n18004_not
g37997 not n18301 ; n18301_not
g37998 not n10435 ; n10435_not
g37999 not n10417 ; n10417_not
g38000 not n10354 ; n10354_not
g38001 not n12046 ; n12046_not
g38002 not n12028 ; n12028_not
g38003 not n20128 ; n20128_not
g38004 not n27022 ; n27022_not
g38005 not n10390 ; n10390_not
g38006 not n20119 ; n20119_not
g38007 not n11722 ; n11722_not
g38008 not n21019 ; n21019_not
g38009 not n12091 ; n12091_not
g38010 not n10408 ; n10408_not
g38011 not n12082 ; n12082_not
g38012 not n11146 ; n11146_not
g38013 not n21190 ; n21190_not
g38014 not n25312 ; n25312_not
g38015 not n11236 ; n11236_not
g38016 not n10912 ; n10912_not
g38017 not n19111 ; n19111_not
g38018 not n17203 ; n17203_not
g38019 not n11227 ; n11227_not
g38020 not n25303 ; n25303_not
g38021 not n11218 ; n11218_not
g38022 not n11209 ; n11209_not
g38023 not n27202 ; n27202_not
g38024 not n12550 ; n12550_not
g38025 not n11182 ; n11182_not
g38026 not n19102 ; n19102_not
g38027 not n11191 ; n11191_not
g38028 not n12604 ; n12604_not
g38029 not n12613 ; n12613_not
g38030 not n18013 ; n18013_not
g38031 not n21208 ; n21208_not
g38032 not n11173 ; n11173_not
g38033 not n10921 ; n10921_not
g38034 not n26221 ; n26221_not
g38035 not n25330 ; n25330_not
g38036 not n20335 ; n20335_not
g38037 not n17230 ; n17230_not
g38038 not n12541 ; n12541_not
g38039 not n11272 ; n11272_not
g38040 not n11281 ; n11281_not
g38041 not n17212 ; n17212_not
g38042 not n19120 ; n19120_not
g38043 not n12253 ; n12253_not
g38044 not n26401 ; n26401_not
g38045 not n17221 ; n17221_not
g38046 not n20236 ; n20236_not
g38047 not n20326 ; n20326_not
g38048 not n27220 ; n27220_not
g38049 not n10903 ; n10903_not
g38050 not n11263 ; n11263_not
g38051 not n11254 ; n11254_not
g38052 not n27211 ; n27211_not
g38053 not n12217 ; n12217_not
g38054 not n25240 ; n25240_not
g38055 not n11056 ; n11056_not
g38056 not n10714 ; n10714_not
g38057 not n17140 ; n17140_not
g38058 not n19012 ; n19012_not
g38059 not n11047 ; n11047_not
g38060 not n11029 ; n11029_not
g38061 not n19003 ; n19003_not
g38062 not n27112 ; n27112_not
g38063 not n20290 ; n20290_not
g38064 not n17005 ; n17005_not
g38065 not n20254 ; n20254_not
g38066 not n25222 ; n25222_not
g38067 not n21244 ; n21244_not
g38068 not n26311 ; n26311_not
g38069 not n20281 ; n20281_not
g38070 not n27121 ; n27121_not
g38071 not n20272 ; n20272_not
g38072 not n26302 ; n26302_not
g38073 not n18121 ; n18121_not
g38074 not n10930 ; n10930_not
g38075 not n12622 ; n12622_not
g38076 not n21217 ; n21217_not
g38077 not n12631 ; n12631_not
g38078 not n18022 ; n18022_not
g38079 not n11155 ; n11155_not
g38080 not n12640 ; n12640_not
g38081 not n18112 ; n18112_not
g38082 not n11137 ; n11137_not
g38083 not n19030 ; n19030_not
g38084 not n11119 ; n11119_not
g38085 not n19021 ; n19021_not
g38086 not n18031 ; n18031_not
g38087 not n11092 ; n11092_not
g38088 not n27103 ; n27103_not
g38089 not n10741 ; n10741_not
g38090 not n11074 ; n11074_not
g38091 not n20245 ; n20245_not
g38092 not n12514 ; n12514_not
g38093 not n12523 ; n12523_not
g38094 not n20218 ; n20218_not
g38095 not n20371 ; n20371_not
g38096 not n21163 ; n21163_not
g38097 not n21172 ; n21172_not
g38098 not n21145 ; n21145_not
g38099 not n11326 ; n11326_not
g38100 not n12532 ; n12532_not
g38101 not n11344 ; n11344_not
g38102 not n26410 ; n26410_not
g38103 not n20353 ; n20353_not
g38104 not n20209 ; n20209_not
g38105 not n20344 ; n20344_not
g38106 not n20362 ; n20362_not
g38107 not n19201 ; n19201_not
g38108 not n11308 ; n11308_not
g38109 not n10634 ; n10634_not
g38110 not n22523 ; n22523_not
g38111 not n10355 ; n10355_not
g38112 not n14036 ; n14036_not
g38113 not n20219 ; n20219_not
g38114 not n11480 ; n11480_not
g38115 not n14441 ; n14441_not
g38116 not n22019 ; n22019_not
g38117 not n18302 ; n18302_not
g38118 not n14252 ; n14252_not
g38119 not n15422 ; n15422_not
g38120 not n26051 ; n26051_not
g38121 not n16007 ; n16007_not
g38122 not n10940 ; n10940_not
g38123 not n23513 ; n23513_not
g38124 not n10643 ; n10643_not
g38125 not n11066 ; n11066_not
g38126 not n16403 ; n16403_not
g38127 not n16016 ; n16016_not
g38128 not n23621 ; n23621_not
g38129 not n14342 ; n14342_not
g38130 not n11417 ; n11417_not
g38131 not n14702 ; n14702_not
g38132 not n22532 ; n22532_not
g38133 not n18311 ; n18311_not
g38134 not n11804 ; n11804_not
g38135 not n16061 ; n16061_not
g38136 not n20192 ; n20192_not
g38137 not n14261 ; n14261_not
g38138 not n23261 ; n23261_not
g38139 not n20660 ; n20660_not
g38140 not n24404 ; n24404_not
g38141 not n26024 ; n26024_not
g38142 not n10625 ; n10625_not
g38143 not n22154 ; n22154_not
g38144 not n11084 ; n11084_not
g38145 not n26033 ; n26033_not
g38146 not n22208 ; n22208_not
g38147 not n16430 ; n16430_not
g38148 not n20642 ; n20642_not
g38149 not n11057 ; n11057_not
g38150 not n16421 ; n16421_not
g38151 not n23504 ; n23504_not
g38152 not n16133 ; n16133_not
g38153 not n10706 ; n10706_not
g38154 not n20606 ; n20606_not
g38155 not n18032 ; n18032_not
g38156 not n26240 ; n26240_not
g38157 not n22505 ; n22505_not
g38158 not n11741 ; n11741_not
g38159 not n14360 ; n14360_not
g38160 not n13721 ; n13721_not
g38161 not n23540 ; n23540_not
g38162 not n10661 ; n10661_not
g38163 not n14225 ; n14225_not
g38164 not n18113 ; n18113_not
g38165 not n10670 ; n10670_not
g38166 not n24071 ; n24071_not
g38167 not n22046 ; n22046_not
g38168 not n14216 ; n14216_not
g38169 not n11408 ; n11408_not
g38170 not n11723 ; n11723_not
g38171 not n20273 ; n20273_not
g38172 not n18050 ; n18050_not
g38173 not n20183 ; n20183_not
g38174 not n14054 ; n14054_not
g38175 not n14081 ; n14081_not
g38176 not n24332 ; n24332_not
g38177 not n18023 ; n18023_not
g38178 not n11138 ; n11138_not
g38179 not n23810 ; n23810_not
g38180 not n22280 ; n22280_not
g38181 not n20570 ; n20570_not
g38182 not n11426 ; n11426_not
g38183 not n11129 ; n11129_not
g38184 not n20624 ; n20624_not
g38185 not n22514 ; n22514_not
g38186 not n11075 ; n11075_not
g38187 not n22028 ; n22028_not
g38188 not n10652 ; n10652_not
g38189 not n24350 ; n24350_not
g38190 not n18041 ; n18041_not
g38191 not n16070 ; n16070_not
g38192 not n23531 ; n23531_not
g38193 not n20453 ; n20453_not
g38194 not n15323 ; n15323_not
g38195 not n16142 ; n16142_not
g38196 not n22037 ; n22037_not
g38197 not n22316 ; n22316_not
g38198 not n24008 ; n24008_not
g38199 not n23900 ; n23900_not
g38200 not n24341 ; n24341_not
g38201 not n11093 ; n11093_not
g38202 not n13370 ; n13370_not
g38203 not n20372 ; n20372_not
g38204 not n11750 ; n11750_not
g38205 not n14351 ; n14351_not
g38206 not n13703 ; n13703_not
g38207 not n20282 ; n20282_not
g38208 not n13550 ; n13550_not
g38209 not n10571 ; n10571_not
g38210 not n23801 ; n23801_not
g38211 not n21821 ; n21821_not
g38212 not n20741 ; n20741_not
g38213 not n26213 ; n26213_not
g38214 not n24314 ; n24314_not
g38215 not n14450 ; n14450_not
g38216 not n21830 ; n21830_not
g38217 not n16034 ; n16034_not
g38218 not n23423 ; n23423_not
g38219 not n16025 ; n16025_not
g38220 not n23432 ; n23432_not
g38221 not n16520 ; n16520_not
g38222 not n10580 ; n10580_not
g38223 not n22613 ; n22613_not
g38224 not n14234 ; n14234_not
g38225 not n20084 ; n20084_not
g38226 not n13460 ; n13460_not
g38227 not n23441 ; n23441_not
g38228 not n18320 ; n18320_not
g38229 not n22604 ; n22604_not
g38230 not n20723 ; n20723_not
g38231 not n16511 ; n16511_not
g38232 not n14315 ; n14315_not
g38233 not n23450 ; n23450_not
g38234 not n14810 ; n14810_not
g38235 not n22640 ; n22640_not
g38236 not n13523 ; n13523_not
g38237 not n22460 ; n22460_not
g38238 not n14801 ; n14801_not
g38239 not n21803 ; n21803_not
g38240 not n17600 ; n17600_not
g38241 not n20066 ; n20066_not
g38242 not n26303 ; n26303_not
g38243 not n24503 ; n24503_not
g38244 not n13640 ; n13640_not
g38245 not n22622 ; n22622_not
g38246 not n10562 ; n10562_not
g38247 not n23405 ; n23405_not
g38248 not n21812 ; n21812_not
g38249 not n20651 ; n20651_not
g38250 not n13532 ; n13532_not
g38251 not n13541 ; n13541_not
g38252 not n10850 ; n10850_not
g38253 not n20750 ; n20750_not
g38254 not n10841 ; n10841_not
g38255 not n22631 ; n22631_not
g38256 not n26312 ; n26312_not
g38257 not n10616 ; n10616_not
g38258 not n24080 ; n24080_not
g38259 not n15701 ; n15701_not
g38260 not n10607 ; n10607_not
g38261 not n16151 ; n16151_not
g38262 not n11831 ; n11831_not
g38263 not n18104 ; n18104_not
g38264 not n21920 ; n21920_not
g38265 not n14720 ; n14720_not
g38266 not n14270 ; n14270_not
g38267 not n22307 ; n22307_not
g38268 not n14333 ; n14333_not
g38269 not n24422 ; n24422_not
g38270 not n22163 ; n22163_not
g38271 not n22541 ; n22541_not
g38272 not n11048 ; n11048_not
g38273 not n20390 ; n20390_not
g38274 not n26015 ; n26015_not
g38275 not n15710 ; n15710_not
g38276 not n23243 ; n23243_not
g38277 not n11822 ; n11822_not
g38278 not n21902 ; n21902_not
g38279 not n13631 ; n13631_not
g38280 not n24440 ; n24440_not
g38281 not n20075 ; n20075_not
g38282 not n16160 ; n16160_not
g38283 not n20381 ; n20381_not
g38284 not n24431 ; n24431_not
g38285 not n14063 ; n14063_not
g38286 not n20714 ; n20714_not
g38287 not n26321 ; n26321_not
g38288 not n20093 ; n20093_not
g38289 not n20705 ; n20705_not
g38290 not n16043 ; n16043_not
g38291 not n13613 ; n13613_not
g38292 not n26006 ; n26006_not
g38293 not n16052 ; n16052_not
g38294 not n26330 ; n26330_not
g38295 not n20291 ; n20291_not
g38296 not n11381 ; n11381_not
g38297 not n21911 ; n21911_not
g38298 not n20255 ; n20255_not
g38299 not n22550 ; n22550_not
g38300 not n14324 ; n14324_not
g38301 not n11264 ; n11264_not
g38302 not n11570 ; n11570_not
g38303 not n20417 ; n20417_not
g38304 not n22091 ; n22091_not
g38305 not n11561 ; n11561_not
g38306 not n20327 ; n20327_not
g38307 not n20237 ; n20237_not
g38308 not n22370 ; n22370_not
g38309 not n26141 ; n26141_not
g38310 not n22127 ; n22127_not
g38311 not n22253 ; n22253_not
g38312 not n24170 ; n24170_not
g38313 not n14540 ; n14540_not
g38314 not n20228 ; n20228_not
g38315 not n11336 ; n11336_not
g38316 not n15602 ; n15602_not
g38317 not n16232 ; n16232_not
g38318 not n22361 ; n22361_not
g38319 not n14135 ; n14135_not
g38320 not n24161 ; n24161_not
g38321 not n11327 ; n11327_not
g38322 not n20471 ; n20471_not
g38323 not n26150 ; n26150_not
g38324 not n13505 ; n13505_not
g38325 not n14531 ; n14531_not
g38326 not n11237 ; n11237_not
g38327 not n24215 ; n24215_not
g38328 not n11246 ; n11246_not
g38329 not n22415 ; n22415_not
g38330 not n20516 ; n20516_not
g38331 not n14153 ; n14153_not
g38332 not n11345 ; n11345_not
g38333 not n16115 ; n16115_not
g38334 not n11255 ; n11255_not
g38335 not n26600 ; n26600_not
g38336 not n20507 ; n20507_not
g38337 not n24044 ; n24044_not
g38338 not n10904 ; n10904_not
g38339 not n18203 ; n18203_not
g38340 not n10751 ; n10751_not
g38341 not n24206 ; n24206_not
g38342 not n26132 ; n26132_not
g38343 not n10526 ; n10526_not
g38344 not n22406 ; n22406_not
g38345 not n13820 ; n13820_not
g38346 not n10463 ; n10463_not
g38347 not n14144 ; n14144_not
g38348 not n20480 ; n20480_not
g38349 not n18131 ; n18131_not
g38350 not n22118 ; n22118_not
g38351 not n22145 ; n22145_not
g38352 not n22064 ; n22064_not
g38353 not n18221 ; n18221_not
g38354 not n20426 ; n20426_not
g38355 not n22352 ; n22352_not
g38356 not n14126 ; n14126_not
g38357 not n24134 ; n24134_not
g38358 not n11309 ; n11309_not
g38359 not n20336 ; n20336_not
g38360 not n16205 ; n16205_not
g38361 not n14504 ; n14504_not
g38362 not n24125 ; n24125_not
g38363 not n18212 ; n18212_not
g38364 not n11525 ; n11525_not
g38365 not n18140 ; n18140_not
g38366 not n11291 ; n11291_not
g38367 not n26222 ; n26222_not
g38368 not n10805 ; n10805_not
g38369 not n22136 ; n22136_not
g38370 not n11516 ; n11516_not
g38371 not n22262 ; n22262_not
g38372 not n22343 ; n22343_not
g38373 not n24116 ; n24116_not
g38374 not n11507 ; n11507_not
g38375 not n23711 ; n23711_not
g38376 not n10436 ; n10436_not
g38377 not n14117 ; n14117_not
g38378 not n23720 ; n23720_not
g38379 not n22172 ; n22172_not
g38380 not n24053 ; n24053_not
g38381 not n11273 ; n11273_not
g38382 not n20174 ; n20174_not
g38383 not n26402 ; n26402_not
g38384 not n11552 ; n11552_not
g38385 not n23702 ; n23702_not
g38386 not n20462 ; n20462_not
g38387 not n10454 ; n10454_not
g38388 not n24152 ; n24152_not
g38389 not n14108 ; n14108_not
g38390 not n14522 ; n14522_not
g38391 not n26231 ; n26231_not
g38392 not n13901 ; n13901_not
g38393 not n16214 ; n16214_not
g38394 not n24143 ; n24143_not
g38395 not n11282 ; n11282_not
g38396 not n14513 ; n14513_not
g38397 not n11543 ; n11543_not
g38398 not n16124 ; n16124_not
g38399 not n22442 ; n22442_not
g38400 not n11444 ; n11444_not
g38401 not n16340 ; n16340_not
g38402 not n26105 ; n26105_not
g38403 not n22073 ; n22073_not
g38404 not n20543 ; n20543_not
g38405 not n11183 ; n11183_not
g38406 not n20129 ; n20129_not
g38407 not n22190 ; n22190_not
g38408 not n14603 ; n14603_not
g38409 not n10922 ; n10922_not
g38410 not n27302 ; n27302_not
g38411 not n18005 ; n18005_not
g38412 not n16322 ; n16322_not
g38413 not n10715 ; n10715_not
g38414 not n11453 ; n11453_not
g38415 not n10724 ; n10724_not
g38416 not n16313 ; n16313_not
g38417 not n24260 ; n24260_not
g38418 not n22226 ; n22226_not
g38419 not n26114 ; n26114_not
g38420 not n24026 ; n24026_not
g38421 not n18122 ; n18122_not
g38422 not n22055 ; n22055_not
g38423 not n11156 ; n11156_not
g38424 not n20246 ; n20246_not
g38425 not n11714 ; n11714_not
g38426 not n14630 ; n14630_not
g38427 not n20561 ; n20561_not
g38428 not n11165 ; n11165_not
g38429 not n10931 ; n10931_not
g38430 not n11705 ; n11705_not
g38431 not n14018 ; n14018_not
g38432 not n14207 ; n14207_not
g38433 not n11435 ; n11435_not
g38434 not n26501 ; n26501_not
g38435 not n14621 ; n14621_not
g38436 not n20552 ; n20552_not
g38437 not n14432 ; n14432_not
g38438 not n20138 ; n20138_not
g38439 not n11174 ; n11174_not
g38440 not n22451 ; n22451_not
g38441 not n24305 ; n24305_not
g38442 not n18014 ; n18014_not
g38443 not n11651 ; n11651_not
g38444 not n11219 ; n11219_not
g38445 not n11462 ; n11462_not
g38446 not n14423 ; n14423_not
g38447 not n11228 ; n11228_not
g38448 not n26042 ; n26042_not
g38449 not n24062 ; n24062_not
g38450 not n11642 ; n11642_not
g38451 not n24233 ; n24233_not
g38452 not n20318 ; n20318_not
g38453 not n26123 ; n26123_not
g38454 not n20525 ; n20525_not
g38455 not n22424 ; n22424_not
g38456 not n20156 ; n20156_not
g38457 not n11633 ; n11633_not
g38458 not n16106 ; n16106_not
g38459 not n11147 ; n11147_not
g38460 not n10913 ; n10913_not
g38461 not n22109 ; n22109_not
g38462 not n11363 ; n11363_not
g38463 not n26510 ; n26510_not
g38464 not n10742 ; n10742_not
g38465 not n14162 ; n14162_not
g38466 not n24224 ; n24224_not
g38467 not n20354 ; n20354_not
g38468 not n26420 ; n26420_not
g38469 not n23630 ; n23630_not
g38470 not n22082 ; n22082_not
g38471 not n11192 ; n11192_not
g38472 not n24251 ; n24251_not
g38473 not n23603 ; n23603_not
g38474 not n14090 ; n14090_not
g38475 not n20408 ; n20408_not
g38476 not n13802 ; n13802_not
g38477 not n15404 ; n15404_not
g38478 not n20534 ; n20534_not
g38479 not n16304 ; n16304_not
g38480 not n20147 ; n20147_not
g38481 not n11660 ; n11660_not
g38482 not n14009 ; n14009_not
g38483 not n22235 ; n22235_not
g38484 not n13811 ; n13811_not
g38485 not n14180 ; n14180_not
g38486 not n23612 ; n23612_not
g38487 not n22334 ; n22334_not
g38488 not n24242 ; n24242_not
g38489 not n12353 ; n12353_not
g38490 not n15080 ; n15080_not
g38491 not n10067 ; n10067_not
g38492 not n22811 ; n22811_not
g38493 not n21425 ; n21425_not
g38494 not n17330 ; n17330_not
g38495 not n19400 ; n19400_not
g38496 not n17321 ; n17321_not
g38497 not n13055 ; n13055_not
g38498 not n23135 ; n23135_not
g38499 not n25421 ; n25421_not
g38500 not n12371 ; n12371_not
g38501 not n10166 ; n10166_not
g38502 not n24800 ; n24800_not
g38503 not n21416 ; n21416_not
g38504 not n10157 ; n10157_not
g38505 not n12380 ; n12380_not
g38506 not n17312 ; n17312_not
g38507 not n10148 ; n10148_not
g38508 not n13037 ; n13037_not
g38509 not n15062 ; n15062_not
g38510 not n12317 ; n12317_not
g38511 not n12326 ; n12326_not
g38512 not n12335 ; n12335_not
g38513 not n10184 ; n10184_not
g38514 not n23144 ; n23144_not
g38515 not n13091 ; n13091_not
g38516 not n21443 ; n21443_not
g38517 not n22910 ; n22910_not
g38518 not n22703 ; n22703_not
g38519 not n13082 ; n13082_not
g38520 not n21434 ; n21434_not
g38521 not n13073 ; n13073_not
g38522 not n21092 ; n21092_not
g38523 not n21371 ; n21371_not
g38524 not n10076 ; n10076_not
g38525 not n12452 ; n12452_not
g38526 not n21380 ; n21380_not
g38527 not n19310 ; n19310_not
g38528 not n15125 ; n15125_not
g38529 not n15350 ; n15350_not
g38530 not n10058 ; n10058_not
g38531 not n10049 ; n10049_not
g38532 not n21362 ; n21362_not
g38533 not n15134 ; n15134_not
g38534 not n12461 ; n12461_not
g38535 not n21128 ; n21128_not
g38536 not n25007 ; n25007_not
g38537 not n12470 ; n12470_not
g38538 not n12290 ; n12290_not
g38539 not n25412 ; n25412_not
g38540 not n10139 ; n10139_not
g38541 not n13028 ; n13028_not
g38542 not n12407 ; n12407_not
g38543 not n15107 ; n15107_not
g38544 not n12416 ; n12416_not
g38545 not n12425 ; n12425_not
g38546 not n12434 ; n12434_not
g38547 not n12731 ; n12731_not
g38548 not n27041 ; n27041_not
g38549 not n25403 ; n25403_not
g38550 not n19031 ; n19031_not
g38551 not n21407 ; n21407_not
g38552 not n10094 ; n10094_not
g38553 not n21119 ; n21119_not
g38554 not n25340 ; n25340_not
g38555 not n12443 ; n12443_not
g38556 not n10085 ; n10085_not
g38557 not n21515 ; n21515_not
g38558 not n21038 ; n21038_not
g38559 not n27032 ; n27032_not
g38560 not n23045 ; n23045_not
g38561 not n23063 ; n23063_not
g38562 not n24710 ; n24710_not
g38563 not n21506 ; n21506_not
g38564 not n17402 ; n17402_not
g38565 not n10292 ; n10292_not
g38566 not n13181 ; n13181_not
g38567 not n12191 ; n12191_not
g38568 not n10283 ; n10283_not
g38569 not n13172 ; n13172_not
g38570 not n12164 ; n12164_not
g38571 not n15008 ; n15008_not
g38572 not n19301 ; n19301_not
g38573 not n15440 ; n15440_not
g38574 not n13226 ; n13226_not
g38575 not n21029 ; n21029_not
g38576 not n12155 ; n12155_not
g38577 not n23180 ; n23180_not
g38578 not n10319 ; n10319_not
g38579 not n13217 ; n13217_not
g38580 not n22901 ; n22901_not
g38581 not n25511 ; n25511_not
g38582 not n13208 ; n13208_not
g38583 not n12173 ; n12173_not
g38584 not n23171 ; n23171_not
g38585 not n12182 ; n12182_not
g38586 not n13190 ; n13190_not
g38587 not n15431 ; n15431_not
g38588 not n17411 ; n17411_not
g38589 not n10238 ; n10238_not
g38590 not n27311 ; n27311_not
g38591 not n15035 ; n15035_not
g38592 not n12254 ; n12254_not
g38593 not n13127 ; n13127_not
g38594 not n12263 ; n12263_not
g38595 not n21056 ; n21056_not
g38596 not n15413 ; n15413_not
g38597 not n12272 ; n12272_not
g38598 not n13118 ; n13118_not
g38599 not n12281 ; n12281_not
g38600 not n18500 ; n18500_not
g38601 not n21065 ; n21065_not
g38602 not n15044 ; n15044_not
g38603 not n13019 ; n13019_not
g38604 not n10193 ; n10193_not
g38605 not n15053 ; n15053_not
g38606 not n10274 ; n10274_not
g38607 not n13163 ; n13163_not
g38608 not n25502 ; n25502_not
g38609 not n12209 ; n12209_not
g38610 not n19112 ; n19112_not
g38611 not n12218 ; n12218_not
g38612 not n13154 ; n13154_not
g38613 not n12227 ; n12227_not
g38614 not n21470 ; n21470_not
g38615 not n17051 ; n17051_not
g38616 not n21461 ; n21461_not
g38617 not n10256 ; n10256_not
g38618 not n13145 ; n13145_not
g38619 not n12236 ; n12236_not
g38620 not n15026 ; n15026_not
g38621 not n13136 ; n13136_not
g38622 not n21047 ; n21047_not
g38623 not n25124 ; n25124_not
g38624 not n15233 ; n15233_not
g38625 not n19040 ; n19040_not
g38626 not n23081 ; n23081_not
g38627 not n12641 ; n12641_not
g38628 not n15242 ; n15242_not
g38629 not n12650 ; n12650_not
g38630 not n21272 ; n21272_not
g38631 not n21227 ; n21227_not
g38632 not n19022 ; n19022_not
g38633 not n15251 ; n15251_not
g38634 not n21263 ; n21263_not
g38635 not n19013 ; n19013_not
g38636 not n15314 ; n15314_not
g38637 not n25160 ; n25160_not
g38638 not n25151 ; n25151_not
g38639 not n27203 ; n27203_not
g38640 not n12830 ; n12830_not
g38641 not n25115 ; n25115_not
g38642 not n19103 ; n19103_not
g38643 not n12605 ; n12605_not
g38644 not n15224 ; n15224_not
g38645 not n12821 ; n12821_not
g38646 not n15215 ; n15215_not
g38647 not n17042 ; n17042_not
g38648 not n12812 ; n12812_not
g38649 not n12542 ; n12542_not
g38650 not n12533 ; n12533_not
g38651 not n12803 ; n12803_not
g38652 not n21209 ; n21209_not
g38653 not n12623 ; n12623_not
g38654 not n25205 ; n25205_not
g38655 not n25223 ; n25223_not
g38656 not n17114 ; n17114_not
g38657 not n23054 ; n23054_not
g38658 not n12722 ; n12722_not
g38659 not n12713 ; n12713_not
g38660 not n27140 ; n27140_not
g38661 not n21245 ; n21245_not
g38662 not n12632 ; n12632_not
g38663 not n27131 ; n27131_not
g38664 not n25214 ; n25214_not
g38665 not n27122 ; n27122_not
g38666 not n17123 ; n17123_not
g38667 not n27113 ; n27113_not
g38668 not n21254 ; n21254_not
g38669 not n15260 ; n15260_not
g38670 not n25241 ; n25241_not
g38671 not n15305 ; n15305_not
g38672 not n27104 ; n27104_not
g38673 not n17006 ; n17006_not
g38674 not n21236 ; n21236_not
g38675 not n23036 ; n23036_not
g38676 not n25034 ; n25034_not
g38677 not n17105 ; n17105_not
g38678 not n12740 ; n12740_not
g38679 not n25232 ; n25232_not
g38680 not n19202 ; n19202_not
g38681 not n21335 ; n21335_not
g38682 not n21164 ; n21164_not
g38683 not n12515 ; n12515_not
g38684 not n23117 ; n23117_not
g38685 not n12614 ; n12614_not
g38686 not n21326 ; n21326_not
g38687 not n15170 ; n15170_not
g38688 not n12920 ; n12920_not
g38689 not n17240 ; n17240_not
g38690 not n21173 ; n21173_not
g38691 not n27230 ; n27230_not
g38692 not n12902 ; n12902_not
g38693 not n17231 ; n17231_not
g38694 not n21137 ; n21137_not
g38695 not n19004 ; n19004_not
g38696 not n25016 ; n25016_not
g38697 not n21353 ; n21353_not
g38698 not n23126 ; n23126_not
g38699 not n21344 ; n21344_not
g38700 not n27050 ; n27050_not
g38701 not n15152 ; n15152_not
g38702 not n19220 ; n19220_not
g38703 not n25025 ; n25025_not
g38704 not n21155 ; n21155_not
g38705 not n23018 ; n23018_not
g38706 not n23090 ; n23090_not
g38707 not n15332 ; n15332_not
g38708 not n21182 ; n21182_not
g38709 not n19121 ; n19121_not
g38710 not n15206 ; n15206_not
g38711 not n25313 ; n25313_not
g38712 not n17015 ; n17015_not
g38713 not n17024 ; n17024_not
g38714 not n17204 ; n17204_not
g38715 not n27212 ; n27212_not
g38716 not n25304 ; n25304_not
g38717 not n17033 ; n17033_not
g38718 not n21191 ; n21191_not
g38719 not n23108 ; n23108_not
g38720 not n21317 ; n21317_not
g38721 not n25043 ; n25043_not
g38722 not n25331 ; n25331_not
g38723 not n25052 ; n25052_not
g38724 not n19130 ; n19130_not
g38725 not n21308 ; n21308_not
g38726 not n25061 ; n25061_not
g38727 not n15341 ; n15341_not
g38728 not n17222 ; n17222_not
g38729 not n25070 ; n25070_not
g38730 not n27221 ; n27221_not
g38731 not n23027 ; n23027_not
g38732 not n17213 ; n17213_not
g38733 not n12560 ; n12560_not
g38734 not n12047 ; n12047_not
g38735 not n12038 ; n12038_not
g38736 not n12029 ; n12029_not
g38737 not n11921 ; n11921_not
g38738 not n10535 ; n10535_not
g38739 not n23342 ; n23342_not
g38740 not n15503 ; n15503_not
g38741 not n13334 ; n13334_not
g38742 not n13325 ; n13325_not
g38743 not n10445 ; n10445_not
g38744 not n11930 ; n11930_not
g38745 not n21614 ; n21614_not
g38746 not n15512 ; n15512_not
g38747 not n21722 ; n21722_not
g38748 not n20930 ; n20930_not
g38749 not n10517 ; n10517_not
g38750 not n21623 ; n21623_not
g38751 not n13451 ; n13451_not
g38752 not n18401 ; n18401_not
g38753 not n12083 ; n12083_not
g38754 not n12092 ; n12092_not
g38755 not n23351 ; n23351_not
g38756 not n21605 ; n21605_not
g38757 not n21740 ; n21740_not
g38758 not n12074 ; n12074_not
g38759 not n12065 ; n12065_not
g38760 not n22433 ; n22433_not
g38761 not n13307 ; n13307_not
g38762 not n22802 ; n22802_not
g38763 not n10418 ; n10418_not
g38764 not n13316 ; n13316_not
g38765 not n21731 ; n21731_not
g38766 not n10427 ; n10427_not
g38767 not n24530 ; n24530_not
g38768 not n23252 ; n23252_not
g38769 not n13424 ; n13424_not
g38770 not n10490 ; n10490_not
g38771 not n24602 ; n24602_not
g38772 not n17510 ; n17510_not
g38773 not n24413 ; n24413_not
g38774 not n16700 ; n16700_not
g38775 not n22730 ; n22730_not
g38776 not n25700 ; n25700_not
g38777 not n23162 ; n23162_not
g38778 not n10481 ; n10481_not
g38779 not n20912 ; n20912_not
g38780 not n13415 ; n13415_not
g38781 not n21650 ; n21650_not
g38782 not n23315 ; n23315_not
g38783 not n27005 ; n27005_not
g38784 not n23306 ; n23306_not
g38785 not n20039 ; n20039_not
g38786 not n13406 ; n13406_not
g38787 not n10472 ; n10472_not
g38788 not n20822 ; n20822_not
g38789 not n22712 ; n22712_not
g38790 not n21713 ; n21713_not
g38791 not n13352 ; n13352_not
g38792 not n10391 ; n10391_not
g38793 not n24620 ; n24620_not
g38794 not n20921 ; n20921_not
g38795 not n13361 ; n13361_not
g38796 not n24611 ; n24611_not
g38797 not n21632 ; n21632_not
g38798 not n15530 ; n15530_not
g38799 not n25610 ; n25610_not
g38800 not n13442 ; n13442_not
g38801 not n20813 ; n20813_not
g38802 not n14900 ; n14900_not
g38803 not n17303 ; n17303_not
g38804 not n13433 ; n13433_not
g38805 not n23324 ; n23324_not
g38806 not n20840 ; n20840_not
g38807 not n21704 ; n21704_not
g38808 not n21641 ; n21641_not
g38809 not n13244 ; n13244_not
g38810 not n23216 ; n23216_not
g38811 not n23360 ; n23360_not
g38812 not n10553 ; n10553_not
g38813 not n16610 ; n16610_not
g38814 not n10382 ; n10382_not
g38815 not n21542 ; n21542_not
g38816 not n24521 ; n24521_not
g38817 not n23225 ; n23225_not
g38818 not n27023 ; n27023_not
g38819 not n21560 ; n21560_not
g38820 not n10364 ; n10364_not
g38821 not n11903 ; n11903_not
g38822 not n21524 ; n21524_not
g38823 not n11912 ; n11912_not
g38824 not n23207 ; n23207_not
g38825 not n12128 ; n12128_not
g38826 not n12119 ; n12119_not
g38827 not n16601 ; n16601_not
g38828 not n13262 ; n13262_not
g38829 not n13253 ; n13253_not
g38830 not n11840 ; n11840_not
g38831 not n24512 ; n24512_not
g38832 not n20057 ; n20057_not
g38833 not n10337 ; n10337_not
g38834 not n10544 ; n10544_not
g38835 not n15611 ; n15611_not
g38836 not n12146 ; n12146_not
g38837 not n23234 ; n23234_not
g38838 not n13235 ; n13235_not
g38839 not n22820 ; n22820_not
g38840 not n13514 ; n13514_not
g38841 not n13280 ; n13280_not
g38842 not n27006 ; n27006_not
g38843 not n23325 ; n23325_not
g38844 not n19140 ; n19140_not
g38845 not n23046 ; n23046_not
g38846 not n22551 ; n22551_not
g38847 not n22722 ; n22722_not
g38848 not n15342 ; n15342_not
g38849 not n22254 ; n22254_not
g38850 not n22542 ; n22542_not
g38851 not n20049 ; n20049_not
g38852 not n16026 ; n16026_not
g38853 not n27123 ; n27123_not
g38854 not n27222 ; n27222_not
g38855 not n23370 ; n23370_not
g38856 not n18312 ; n18312_not
g38857 not n10950 ; n10950_not
g38858 not n18132 ; n18132_not
g38859 not n23037 ; n23037_not
g38860 not n22632 ; n22632_not
g38861 not n22560 ; n22560_not
g38862 not n23811 ; n23811_not
g38863 not n15207 ; n15207_not
g38864 not n10473 ; n10473_not
g38865 not n23604 ; n23604_not
g38866 not n15630 ; n15630_not
g38867 not n22713 ; n22713_not
g38868 not n22461 ; n22461_not
g38869 not n19113 ; n19113_not
g38870 not n18150 ; n18150_not
g38871 not n20256 ; n20256_not
g38872 not n14325 ; n14325_not
g38873 not n26322 ; n26322_not
g38874 not n22641 ; n22641_not
g38875 not n18600 ; n18600_not
g38876 not n15333 ; n15333_not
g38877 not n23109 ; n23109_not
g38878 not n14406 ; n14406_not
g38879 not n15702 ; n15702_not
g38880 not n10482 ; n10482_not
g38881 not n10356 ; n10356_not
g38882 not n23316 ; n23316_not
g38883 not n26403 ; n26403_not
g38884 not n20265 ; n20265_not
g38885 not n15612 ; n15612_not
g38886 not n18051 ; n18051_not
g38887 not n27132 ; n27132_not
g38888 not n18141 ; n18141_not
g38889 not n27060 ; n27060_not
g38890 not n14721 ; n14721_not
g38891 not n26313 ; n26313_not
g38892 not n22263 ; n22263_not
g38893 not n20229 ; n20229_not
g38894 not n23055 ; n23055_not
g38895 not n23802 ; n23802_not
g38896 not n27231 ; n27231_not
g38897 not n19122 ; n19122_not
g38898 not n14811 ; n14811_not
g38899 not n27114 ; n27114_not
g38900 not n14316 ; n14316_not
g38901 not n11436 ; n11436_not
g38902 not n15603 ; n15603_not
g38903 not n10554 ; n10554_not
g38904 not n19131 ; n19131_not
g38905 not n15180 ; n15180_not
g38906 not n10491 ; n10491_not
g38907 not n15621 ; n15621_not
g38908 not n20247 ; n20247_not
g38909 not n10545 ; n10545_not
g38910 not n27150 ; n27150_not
g38911 not n10581 ; n10581_not
g38912 not n19032 ; n19032_not
g38913 not n20058 ; n20058_not
g38914 not n10536 ; n10536_not
g38915 not n15306 ; n15306_not
g38916 not n19041 ; n19041_not
g38917 not n15234 ; n15234_not
g38918 not n23901 ; n23901_not
g38919 not n10932 ; n10932_not
g38920 not n22614 ; n22614_not
g38921 not n10563 ; n10563_not
g38922 not n15261 ; n15261_not
g38923 not n10941 ; n10941_not
g38924 not n18330 ; n18330_not
g38925 not n10923 ; n10923_not
g38926 not n14370 ; n14370_not
g38927 not n15054 ; n15054_not
g38928 not n26340 ; n26340_not
g38929 not n14343 ; n14343_not
g38930 not n23343 ; n23343_not
g38931 not n15252 ; n15252_not
g38932 not n23703 ; n23703_not
g38933 not n19014 ; n19014_not
g38934 not n22227 ; n22227_not
g38935 not n22623 ; n22623_not
g38936 not n16008 ; n16008_not
g38937 not n10572 ; n10572_not
g38938 not n14361 ; n14361_not
g38939 not n14352 ; n14352_not
g38940 not n19023 ; n19023_not
g38941 not n20076 ; n20076_not
g38942 not n22650 ; n22650_not
g38943 not n27042 ; n27042_not
g38944 not n18114 ; n18114_not
g38945 not n23424 ; n23424_not
g38946 not n23352 ; n23352_not
g38947 not n10752 ; n10752_not
g38948 not n15243 ; n15243_not
g38949 not n14901 ; n14901_not
g38950 not n27033 ; n27033_not
g38951 not n22236 ; n22236_not
g38952 not n19005 ; n19005_not
g38953 not n23442 ; n23442_not
g38954 not n22380 ; n22380_not
g38955 not n14334 ; n14334_not
g38956 not n23361 ; n23361_not
g38957 not n27141 ; n27141_not
g38958 not n27204 ; n27204_not
g38959 not n23082 ; n23082_not
g38960 not n20067 ; n20067_not
g38961 not n10914 ; n10914_not
g38962 not n20238 ; n20238_not
g38963 not n14820 ; n14820_not
g38964 not n23820 ; n23820_not
g38965 not n27213 ; n27213_not
g38966 not n23433 ; n23433_not
g38967 not n26331 ; n26331_not
g38968 not n23460 ; n23460_not
g38969 not n10509 ; n10509_not
g38970 not n18105 ; n18105_not
g38971 not n20085 ; n20085_not
g38972 not n14730 ; n14730_not
g38973 not n23064 ; n23064_not
g38974 not n23406 ; n23406_not
g38975 not n15270 ; n15270_not
g38976 not n19050 ; n19050_not
g38977 not n22605 ; n22605_not
g38978 not n18123 ; n18123_not
g38979 not n15324 ; n15324_not
g38980 not n18321 ; n18321_not
g38981 not n15225 ; n15225_not
g38982 not n16017 ; n16017_not
g38983 not n23451 ; n23451_not
g38984 not n10518 ; n10518_not
g38985 not n15216 ; n15216_not
g38986 not n14541 ; n14541_not
g38987 not n22308 ; n22308_not
g38988 not n22812 ; n22812_not
g38989 not n15414 ; n15414_not
g38990 not n22371 ; n22371_not
g38991 not n15036 ; n15036_not
g38992 not n18402 ; n18402_not
g38993 not n10680 ; n10680_not
g38994 not n27312 ; n27312_not
g38995 not n22821 ; n22821_not
g38996 not n10770 ; n10770_not
g38997 not n14550 ; n14550_not
g38998 not n10239 ; n10239_not
g38999 not n20166 ; n20166_not
g39000 not n18240 ; n18240_not
g39001 not n10248 ; n10248_not
g39002 not n22911 ; n22911_not
g39003 not n15027 ; n15027_not
g39004 not n14631 ; n14631_not
g39005 not n22830 ; n22830_not
g39006 not n10329 ; n10329_not
g39007 not n23226 ; n23226_not
g39008 not n15711 ; n15711_not
g39009 not n10383 ; n10383_not
g39010 not n23640 ; n23640_not
g39011 not n10257 ; n10257_not
g39012 not n22920 ; n22920_not
g39013 not n18222 ; n18222_not
g39014 not n19410 ; n19410_not
g39015 not n15072 ; n15072_not
g39016 not n18213 ; n18213_not
g39017 not n14514 ; n14514_not
g39018 not n22353 ; n22353_not
g39019 not n10419 ; n10419_not
g39020 not n22803 ; n22803_not
g39021 not n10185 ; n10185_not
g39022 not n15063 ; n15063_not
g39023 not n14523 ; n14523_not
g39024 not n23541 ; n23541_not
g39025 not n23550 ; n23550_not
g39026 not n20175 ; n20175_not
g39027 not n18510 ; n18510_not
g39028 not n18231 ; n18231_not
g39029 not n10194 ; n10194_not
g39030 not n10662 ; n10662_not
g39031 not n18501 ; n18501_not
g39032 not n23244 ; n23244_not
g39033 not n14532 ; n14532_not
g39034 not n10671 ; n10671_not
g39035 not n14640 ; n14640_not
g39036 not n15045 ; n15045_not
g39037 not n22362 ; n22362_not
g39038 not n15810 ; n15810_not
g39039 not n22425 ; n22425_not
g39040 not n26610 ; n26610_not
g39041 not n10293 ; n10293_not
g39042 not n20139 ; n20139_not
g39043 not n23208 ; n23208_not
g39044 not n14613 ; n14613_not
g39045 not n10176 ; n10176_not
g39046 not n15450 ; n15450_not
g39047 not n14604 ; n14604_not
g39048 not n23172 ; n23172_not
g39049 not n15432 ; n15432_not
g39050 not n15423 ; n15423_not
g39051 not n10707 ; n10707_not
g39052 not n10338 ; n10338_not
g39053 not n23019 ; n23019_not
g39054 not n23190 ; n23190_not
g39055 not n20148 ; n20148_not
g39056 not n10725 ; n10725_not
g39057 not n23181 ; n23181_not
g39058 not n22704 ; n22704_not
g39059 not n10158 ; n10158_not
g39060 not n18411 ; n18411_not
g39061 not n23217 ; n23217_not
g39062 not n22416 ; n22416_not
g39063 not n10275 ; n10275_not
g39064 not n26601 ; n26601_not
g39065 not n23631 ; n23631_not
g39066 not n10374 ; n10374_not
g39067 not n23622 ; n23622_not
g39068 not n20157 ; n20157_not
g39069 not n15009 ; n15009_not
g39070 not n27024 ; n27024_not
g39071 not n22452 ; n22452_not
g39072 not n10365 ; n10365_not
g39073 not n10743 ; n10743_not
g39074 not n10284 ; n10284_not
g39075 not n22434 ; n22434_not
g39076 not n19311 ; n19311_not
g39077 not n15801 ; n15801_not
g39078 not n22443 ; n22443_not
g39079 not n15144 ; n15144_not
g39080 not n23127 ; n23127_not
g39081 not n26502 ; n26502_not
g39082 not n10842 ; n10842_not
g39083 not n10455 ; n10455_not
g39084 not n15540 ; n15540_not
g39085 not n14451 ; n14451_not
g39086 not n15720 ; n15720_not
g39087 not n19302 ; n19302_not
g39088 not n15351 ; n15351_not
g39089 not n15135 ; n15135_not
g39090 not n15081 ; n15081_not
g39091 not n23280 ; n23280_not
g39092 not n22290 ; n22290_not
g39093 not n15360 ; n15360_not
g39094 not n20193 ; n20193_not
g39095 not n14460 ; n14460_not
g39096 not n10626 ; n10626_not
g39097 not n23505 ; n23505_not
g39098 not n15531 ; n15531_not
g39099 not n27303 ; n27303_not
g39100 not n15126 ; n15126_not
g39101 not n22317 ; n22317_not
g39102 not n26421 ; n26421_not
g39103 not n15171 ; n15171_not
g39104 not n14424 ; n14424_not
g39105 not n23307 ; n23307_not
g39106 not n22038 ; n22038_not
g39107 not n22272 ; n22272_not
g39108 not n10464 ; n10464_not
g39109 not n27051 ; n27051_not
g39110 not n27240 ; n27240_not
g39111 not n26430 ; n26430_not
g39112 not n19203 ; n19203_not
g39113 not n14703 ; n14703_not
g39114 not n22281 ; n22281_not
g39115 not n10860 ; n10860_not
g39116 not n19212 ; n19212_not
g39117 not n15153 ; n15153_not
g39118 not n10617 ; n10617_not
g39119 not n19221 ; n19221_not
g39120 not n22533 ; n22533_not
g39121 not n14442 ; n14442_not
g39122 not n27015 ; n27015_not
g39123 not n19230 ; n19230_not
g39124 not n22731 ; n22731_not
g39125 not n22524 ; n22524_not
g39126 not n23721 ; n23721_not
g39127 not n15513 ; n15513_not
g39128 not n10149 ; n10149_not
g39129 not n10392 ; n10392_not
g39130 not n18204 ; n18204_not
g39131 not n10815 ; n10815_not
g39132 not n23523 ; n23523_not
g39133 not n10446 ; n10446_not
g39134 not n10806 ; n10806_not
g39135 not n15504 ; n15504_not
g39136 not n23712 ; n23712_not
g39137 not n23136 ; n23136_not
g39138 not n15090 ; n15090_not
g39139 not n19401 ; n19401_not
g39140 not n26511 ; n26511_not
g39141 not n10437 ; n10437_not
g39142 not n10653 ; n10653_not
g39143 not n23532 ; n23532_not
g39144 not n14505 ; n14505_not
g39145 not n22344 ; n22344_not
g39146 not n20094 ; n20094_not
g39147 not n22506 ; n22506_not
g39148 not n10068 ; n10068_not
g39149 not n10077 ; n10077_not
g39150 not n10086 ; n10086_not
g39151 not n22326 ; n22326_not
g39152 not n10824 ; n10824_not
g39153 not n22740 ; n22740_not
g39154 not n10635 ; n10635_not
g39155 not n15117 ; n15117_not
g39156 not n19320 ; n19320_not
g39157 not n23514 ; n23514_not
g39158 not n23163 ; n23163_not
g39159 not n14910 ; n14910_not
g39160 not n23262 ; n23262_not
g39161 not n15108 ; n15108_not
g39162 not n22335 ; n22335_not
g39163 not n14118 ; n14118_not
g39164 not n10644 ; n10644_not
g39165 not n23730 ; n23730_not
g39166 not n15900 ; n15900_not
g39167 not n14217 ; n14217_not
g39168 not n20913 ; n20913_not
g39169 not n17511 ; n17511_not
g39170 not n25620 ; n25620_not
g39171 not n21642 ; n21642_not
g39172 not n16701 ; n16701_not
g39173 not n13380 ; n13380_not
g39174 not n25611 ; n25611_not
g39175 not n16710 ; n16710_not
g39176 not n13371 ; n13371_not
g39177 not n21633 ; n21633_not
g39178 not n25602 ; n25602_not
g39179 not n17502 ; n17502_not
g39180 not n21624 ; n21624_not
g39181 not n20922 ; n20922_not
g39182 not n24621 ; n24621_not
g39183 not n13353 ; n13353_not
g39184 not n25305 ; n25305_not
g39185 not n20931 ; n20931_not
g39186 not n20940 ; n20940_not
g39187 not n21615 ; n21615_not
g39188 not n13335 ; n13335_not
g39189 not n20724 ; n20724_not
g39190 not n25530 ; n25530_not
g39191 not n13326 ; n13326_not
g39192 not n17232 ; n17232_not
g39193 not n11922 ; n11922_not
g39194 not n24540 ; n24540_not
g39195 not n21507 ; n21507_not
g39196 not n11931 ; n11931_not
g39197 not n13452 ; n13452_not
g39198 not n20823 ; n20823_not
g39199 not n25710 ; n25710_not
g39200 not n21714 ; n21714_not
g39201 not n13443 ; n13443_not
g39202 not n13227 ; n13227_not
g39203 not n21705 ; n21705_not
g39204 not n11940 ; n11940_not
g39205 not n20841 ; n20841_not
g39206 not n13425 ; n13425_not
g39207 not n20850 ; n20850_not
g39208 not n25701 ; n25701_not
g39209 not n11580 ; n11580_not
g39210 not n13281 ; n13281_not
g39211 not n20742 ; n20742_not
g39212 not n13407 ; n13407_not
g39213 not n17520 ; n17520_not
g39214 not n21651 ; n21651_not
g39215 not n13263 ; n13263_not
g39216 not n16800 ; n16800_not
g39217 not n21525 ; n21525_not
g39218 not n13254 ; n13254_not
g39219 not n12129 ; n12129_not
g39220 not n13245 ; n13245_not
g39221 not n25521 ; n25521_not
g39222 not n12138 ; n12138_not
g39223 not n17430 ; n17430_not
g39224 not n25512 ; n25512_not
g39225 not n13236 ; n13236_not
g39226 not n12147 ; n12147_not
g39227 not n21516 ; n21516_not
g39228 not n17421 ; n17421_not
g39229 not n13209 ; n13209_not
g39230 not n13218 ; n13218_not
g39231 not n12165 ; n12165_not
g39232 not n17412 ; n17412_not
g39233 not n12174 ; n12174_not
g39234 not n12048 ; n12048_not
g39235 not n13308 ; n13308_not
g39236 not n13317 ; n13317_not
g39237 not n12039 ; n12039_not
g39238 not n12057 ; n12057_not
g39239 not n21606 ; n21606_not
g39240 not n20751 ; n20751_not
g39241 not n12066 ; n12066_not
g39242 not n12075 ; n12075_not
g39243 not n24630 ; n24630_not
g39244 not n12084 ; n12084_not
g39245 not n12093 ; n12093_not
g39246 not n21471 ; n21471_not
g39247 not n13290 ; n13290_not
g39248 not n21570 ; n21570_not
g39249 not n21561 ; n21561_not
g39250 not n21552 ; n21552_not
g39251 not n11841 ; n11841_not
g39252 not n21543 ; n21543_not
g39253 not n13272 ; n13272_not
g39254 not n21534 ; n21534_not
g39255 not n20355 ; n20355_not
g39256 not n11823 ; n11823_not
g39257 not n21912 ; n21912_not
g39258 not n21660 ; n21660_not
g39259 not n13614 ; n13614_not
g39260 not n13164 ; n13164_not
g39261 not n26007 ; n26007_not
g39262 not n21903 ; n21903_not
g39263 not n13605 ; n13605_not
g39264 not n24423 ; n24423_not
g39265 not n11850 ; n11850_not
g39266 not n24351 ; n24351_not
g39267 not n20715 ; n20715_not
g39268 not n11670 ; n11670_not
g39269 not n24432 ; n24432_not
g39270 not n16503 ; n16503_not
g39271 not n24441 ; n24441_not
g39272 not n24450 ; n24450_not
g39273 not n16512 ; n16512_not
g39274 not n16143 ; n16143_not
g39275 not n20445 ; n20445_not
g39276 not n24360 ; n24360_not
g39277 not n16404 ; n16404_not
g39278 not n24243 ; n24243_not
g39279 not n26052 ; n26052_not
g39280 not n20634 ; n20634_not
g39281 not n13434 ; n13434_not
g39282 not n16422 ; n16422_not
g39283 not n17700 ; n17700_not
g39284 not n20643 ; n20643_not
g39285 not n20409 ; n20409_not
g39286 not n26025 ; n26025_not
g39287 not n24405 ; n24405_not
g39288 not n11454 ; n11454_not
g39289 not n16440 ; n16440_not
g39290 not n13650 ; n13650_not
g39291 not n20661 ; n20661_not
g39292 not n13641 ; n13641_not
g39293 not n26016 ; n26016_not
g39294 not n21732 ; n21732_not
g39295 not n21813 ; n21813_not
g39296 not n16305 ; n16305_not
g39297 not n13632 ; n13632_not
g39298 not n21723 ; n21723_not
g39299 not n11553 ; n11553_not
g39300 not n13515 ; n13515_not
g39301 not n25800 ; n25800_not
g39302 not n21750 ; n21750_not
g39303 not n13506 ; n13506_not
g39304 not n11904 ; n11904_not
g39305 not n20805 ; n20805_not
g39306 not n24513 ; n24513_not
g39307 not n16602 ; n16602_not
g39308 not n20814 ; n20814_not
g39309 not n24522 ; n24522_not
g39310 not n16611 ; n16611_not
g39311 not n21741 ; n21741_not
g39312 not n13092 ; n13092_not
g39313 not n13470 ; n13470_not
g39314 not n24414 ; n24414_not
g39315 not n24531 ; n24531_not
g39316 not n20553 ; n20553_not
g39317 not n16521 ; n16521_not
g39318 not n13461 ; n13461_not
g39319 not n20733 ; n20733_not
g39320 not n16530 ; n16530_not
g39321 not n21840 ; n21840_not
g39322 not n21831 ; n21831_not
g39323 not n13560 ; n13560_not
g39324 not n21822 ; n21822_not
g39325 not n13551 ; n13551_not
g39326 not n17610 ; n17610_not
g39327 not n20652 ; n20652_not
g39328 not n13542 ; n13542_not
g39329 not n11562 ; n11562_not
g39330 not n13533 ; n13533_not
g39331 not n21804 ; n21804_not
g39332 not n17601 ; n17601_not
g39333 not n24504 ; n24504_not
g39334 not n20760 ; n20760_not
g39335 not n13524 ; n13524_not
g39336 not n20616 ; n20616_not
g39337 not n12264 ; n12264_not
g39338 not n25062 ; n25062_not
g39339 not n17223 ; n17223_not
g39340 not n25071 ; n25071_not
g39341 not n12552 ; n12552_not
g39342 not n25323 ; n25323_not
g39343 not n25080 ; n25080_not
g39344 not n12561 ; n12561_not
g39345 not n17214 ; n17214_not
g39346 not n21183 ; n21183_not
g39347 not n17007 ; n17007_not
g39348 not n12228 ; n12228_not
g39349 not n25314 ; n25314_not
g39350 not n12570 ; n12570_not
g39351 not n17016 ; n17016_not
g39352 not n17205 ; n17205_not
g39353 not n17025 ; n17025_not
g39354 not n12840 ; n12840_not
g39355 not n12831 ; n12831_not
g39356 not n21192 ; n21192_not
g39357 not n12480 ; n12480_not
g39358 not n25017 ; n25017_not
g39359 not n21354 ; n21354_not
g39360 not n21345 ; n21345_not
g39361 not n25350 ; n25350_not
g39362 not n17250 ; n17250_not
g39363 not n21336 ; n21336_not
g39364 not n12507 ; n12507_not
g39365 not n12930 ; n12930_not
g39366 not n12516 ; n12516_not
g39367 not n21165 ; n21165_not
g39368 not n21327 ; n21327_not
g39369 not n12921 ; n12921_not
g39370 not n12615 ; n12615_not
g39371 not n12912 ; n12912_not
g39372 not n25035 ; n25035_not
g39373 not n12534 ; n12534_not
g39374 not n12903 ; n12903_not
g39375 not n21318 ; n21318_not
g39376 not n25044 ; n25044_not
g39377 not n25332 ; n25332_not
g39378 not n25053 ; n25053_not
g39379 not n25251 ; n25251_not
g39380 not n21255 ; n21255_not
g39381 not n25143 ; n25143_not
g39382 not n25170 ; n25170_not
g39383 not n17160 ; n17160_not
g39384 not n12660 ; n12660_not
g39385 not n25242 ; n25242_not
g39386 not n12750 ; n12750_not
g39387 not n12354 ; n12354_not
g39388 not n25233 ; n25233_not
g39389 not n12741 ; n12741_not
g39390 not n17142 ; n17142_not
g39391 not n17106 ; n17106_not
g39392 not n12732 ; n12732_not
g39393 not n25224 ; n25224_not
g39394 not n17115 ; n17115_not
g39395 not n17133 ; n17133_not
g39396 not n17124 ; n17124_not
g39397 not n21246 ; n21246_not
g39398 not n25215 ; n25215_not
g39399 not n25116 ; n25116_not
g39400 not n21291 ; n21291_not
g39401 not n12822 ; n12822_not
g39402 not n12606 ; n12606_not
g39403 not n17043 ; n17043_not
g39404 not n12813 ; n12813_not
g39405 not n12453 ; n12453_not
g39406 not n17052 ; n17052_not
g39407 not n12804 ; n12804_not
g39408 not n12624 ; n12624_not
g39409 not n25125 ; n25125_not
g39410 not n25260 ; n25260_not
g39411 not n21282 ; n21282_not
g39412 not n12633 ; n12633_not
g39413 not n12642 ; n12642_not
g39414 not n25134 ; n25134_not
g39415 not n21273 ; n21273_not
g39416 not n17070 ; n17070_not
g39417 not n21228 ; n21228_not
g39418 not n12417 ; n12417_not
g39419 not n21264 ; n21264_not
g39420 not n25152 ; n25152_not
g39421 not n25161 ; n25161_not
g39422 not n12237 ; n12237_not
g39423 not n13137 ; n13137_not
g39424 not n21462 ; n21462_not
g39425 not n21048 ; n21048_not
g39426 not n13128 ; n13128_not
g39427 not n12255 ; n12255_not
g39428 not n25404 ; n25404_not
g39429 not n21057 ; n21057_not
g39430 not n12273 ; n12273_not
g39431 not n13119 ; n13119_not
g39432 not n12282 ; n12282_not
g39433 not n21066 ; n21066_not
g39434 not n12291 ; n12291_not
g39435 not n21075 ; n21075_not
g39436 not n25440 ; n25440_not
g39437 not n12318 ; n12318_not
g39438 not n21453 ; n21453_not
g39439 not n12336 ; n12336_not
g39440 not n12183 ; n12183_not
g39441 not n13191 ; n13191_not
g39442 not n21039 ; n21039_not
g39443 not n17403 ; n17403_not
g39444 not n13182 ; n13182_not
g39445 not n25503 ; n25503_not
g39446 not n24711 ; n24711_not
g39447 not n11814 ; n11814_not
g39448 not n12192 ; n12192_not
g39449 not n13173 ; n13173_not
g39450 not n21480 ; n21480_not
g39451 not n12219 ; n12219_not
g39452 not n24720 ; n24720_not
g39453 not n13155 ; n13155_not
g39454 not n13146 ; n13146_not
g39455 not n12435 ; n12435_not
g39456 not n24810 ; n24810_not
g39457 not n21408 ; n21408_not
g39458 not n12444 ; n12444_not
g39459 not n21390 ; n21390_not
g39460 not n21381 ; n21381_not
g39461 not n24900 ; n24900_not
g39462 not n21372 ; n21372_not
g39463 not n21363 ; n21363_not
g39464 not n25341 ; n25341_not
g39465 not n12462 ; n12462_not
g39466 not n25008 ; n25008_not
g39467 not n12471 ; n12471_not
g39468 not n21138 ; n21138_not
g39469 not n21444 ; n21444_not
g39470 not n21084 ; n21084_not
g39471 not n21435 ; n21435_not
g39472 not n21093 ; n21093_not
g39473 not n17331 ; n17331_not
g39474 not n21426 ; n21426_not
g39475 not n17322 ; n17322_not
g39476 not n13056 ; n13056_not
g39477 not n25422 ; n25422_not
g39478 not n12381 ; n12381_not
g39479 not n21417 ; n21417_not
g39480 not n17313 ; n17313_not
g39481 not n13038 ; n13038_not
g39482 not n12390 ; n12390_not
g39483 not n17304 ; n17304_not
g39484 not n13029 ; n13029_not
g39485 not n12327 ; n12327_not
g39486 not n26205 ; n26205_not
g39487 not n11391 ; n11391_not
g39488 not n11445 ; n11445_not
g39489 not n11463 ; n11463_not
g39490 not n24090 ; n24090_not
g39491 not n22146 ; n22146_not
g39492 not n20418 ; n20418_not
g39493 not n24054 ; n24054_not
g39494 not n11364 ; n11364_not
g39495 not n11229 ; n11229_not
g39496 not n26070 ; n26070_not
g39497 not n11490 ; n11490_not
g39498 not n20427 ; n20427_not
g39499 not n24108 ; n24108_not
g39500 not n20436 ; n20436_not
g39501 not n24117 ; n24117_not
g39502 not n11517 ; n11517_not
g39503 not n16152 ; n16152_not
g39504 not n14064 ; n14064_not
g39505 not n20373 ; n20373_not
g39506 not n24081 ; n24081_not
g39507 not n26214 ; n26214_not
g39508 not n22164 ; n22164_not
g39509 not n14055 ; n14055_not
g39510 not n16161 ; n16161_not
g39511 not n20382 ; n20382_not
g39512 not n22155 ; n22155_not
g39513 not n20391 ; n20391_not
g39514 not n14037 ; n14037_not
g39515 not n11409 ; n11409_not
g39516 not n11418 ; n11418_not
g39517 not n16170 ; n16170_not
g39518 not n14028 ; n14028_not
g39519 not n11427 ; n11427_not
g39520 not n14019 ; n14019_not
g39521 not n22128 ; n22128_not
g39522 not n24171 ; n24171_not
g39523 not n16242 ; n16242_not
g39524 not n20472 ; n20472_not
g39525 not n26142 ; n26142_not
g39526 not n11571 ; n11571_not
g39527 not n16251 ; n16251_not
g39528 not n22119 ; n22119_not
g39529 not n20481 ; n20481_not
g39530 not n20490 ; n20490_not
g39531 not n26133 ; n26133_not
g39532 not n20274 ; n20274_not
g39533 not n24207 ; n24207_not
g39534 not n16260 ; n16260_not
g39535 not n26124 ; n26124_not
g39536 not n11607 ; n11607_not
g39537 not n11616 ; n11616_not
g39538 not n24225 ; n24225_not
g39539 not n20328 ; n20328_not
g39540 not n24135 ; n24135_not
g39541 not n16206 ; n16206_not
g39542 not n11535 ; n11535_not
g39543 not n20454 ; n20454_not
g39544 not n26160 ; n26160_not
g39545 not n22137 ; n22137_not
g39546 not n11544 ; n11544_not
g39547 not n24144 ; n24144_not
g39548 not n16215 ; n16215_not
g39549 not n13902 ; n13902_not
g39550 not n11508 ; n11508_not
g39551 not n24153 ; n24153_not
g39552 not n16224 ; n16224_not
g39553 not n13920 ; n13920_not
g39554 not n24162 ; n24162_not
g39555 not n16233 ; n16233_not
g39556 not n18042 ; n18042_not
g39557 not n11085 ; n11085_not
g39558 not n16071 ; n16071_not
g39559 not n11094 ; n11094_not
g39560 not n24009 ; n24009_not
g39561 not n18033 ; n18033_not
g39562 not n14226 ; n14226_not
g39563 not n26250 ; n26250_not
g39564 not n26241 ; n26241_not
g39565 not n11148 ; n11148_not
g39566 not n16080 ; n16080_not
g39567 not n11157 ; n11157_not
g39568 not n11166 ; n11166_not
g39569 not n14208 ; n14208_not
g39570 not n22191 ; n22191_not
g39571 not n18015 ; n18015_not
g39572 not n11184 ; n11184_not
g39573 not n14190 ; n14190_not
g39574 not n18006 ; n18006_not
g39575 not n24018 ; n24018_not
g39576 not n14307 ; n14307_not
g39577 not n16035 ; n16035_not
g39578 not n14235 ; n14235_not
g39579 not n22218 ; n22218_not
g39580 not n20283 ; n20283_not
g39581 not n16044 ; n16044_not
g39582 not n18060 ; n18060_not
g39583 not n20292 ; n20292_not
g39584 not n14280 ; n14280_not
g39585 not n16053 ; n16053_not
g39586 not n14271 ; n14271_not
g39587 not n16062 ; n16062_not
g39588 not n10716 ; n10716_not
g39589 not n11049 ; n11049_not
g39590 not n22209 ; n22209_not
g39591 not n11058 ; n11058_not
g39592 not n14253 ; n14253_not
g39593 not n11067 ; n11067_not
g39594 not n14127 ; n14127_not
g39595 not n20337 ; n20337_not
g39596 not n26223 ; n26223_not
g39597 not n11292 ; n11292_not
g39598 not n11319 ; n11319_not
g39599 not n14109 ; n14109_not
g39600 not n11328 ; n11328_not
g39601 not n11337 ; n11337_not
g39602 not n11346 ; n11346_not
g39603 not n11355 ; n11355_not
g39604 not n24063 ; n24063_not
g39605 not n26043 ; n26043_not
g39606 not n16134 ; n16134_not
g39607 not n14082 ; n14082_not
g39608 not n11373 ; n11373_not
g39609 not n24072 ; n24072_not
g39610 not n26151 ; n26151_not
g39611 not n24027 ; n24027_not
g39612 not n22182 ; n22182_not
g39613 not n14181 ; n14181_not
g39614 not n20319 ; n20319_not
g39615 not n24036 ; n24036_not
g39616 not n16107 ; n16107_not
g39617 not n14163 ; n14163_not
g39618 not n11238 ; n11238_not
g39619 not n11247 ; n11247_not
g39620 not n14154 ; n14154_not
g39621 not n11256 ; n11256_not
g39622 not n24045 ; n24045_not
g39623 not n14145 ; n14145_not
g39624 not n11265 ; n11265_not
g39625 not n13821 ; n13821_not
g39626 not n26232 ; n26232_not
g39627 not n11274 ; n11274_not
g39628 not n14136 ; n14136_not
g39629 not n11283 ; n11283_not
g39630 not n16125 ; n16125_not
g39631 not n24315 ; n24315_not
g39632 not n20607 ; n20607_not
g39633 not n16341 ; n16341_not
g39634 not n22029 ; n22029_not
g39635 not n13803 ; n13803_not
g39636 not n26106 ; n26106_not
g39637 not n16314 ; n16314_not
g39638 not n11742 ; n11742_not
g39639 not n11724 ; n11724_not
g39640 not n11733 ; n11733_not
g39641 not n11760 ; n11760_not
g39642 not n22092 ; n22092_not
g39643 not n11751 ; n11751_not
g39644 not n13722 ; n13722_not
g39645 not n26115 ; n26115_not
g39646 not n24270 ; n24270_not
g39647 not n13812 ; n13812_not
g39648 not n13713 ; n13713_not
g39649 not n22056 ; n22056_not
g39650 not n11661 ; n11661_not
g39651 not n22074 ; n22074_not
g39652 not n11652 ; n11652_not
g39653 not n20562 ; n20562_not
g39654 not n13704 ; n13704_not
g39655 not n16332 ; n16332_not
g39656 not n13740 ; n13740_not
g39657 not n11715 ; n11715_not
g39658 not n20535 ; n20535_not
g39659 not n11706 ; n11706_not
g39660 not n26061 ; n26061_not
g39661 not n20526 ; n20526_not
g39662 not n11634 ; n11634_not
g39663 not n24252 ; n24252_not
g39664 not n24306 ; n24306_not
g39665 not n24333 ; n24333_not
g39666 not n20580 ; n20580_not
g39667 not n13830 ; n13830_not
g39668 not n22047 ; n22047_not
g39669 not n20571 ; n20571_not
g39670 not n20544 ; n20544_not
g39671 not n16323 ; n16323_not
g39672 not n24234 ; n24234_not
g39673 not n11481 ; n11481_not
g39674 not n20625 ; n20625_not
g39675 not n21355 ; n21355_not
g39676 not n16108 ; n16108_not
g39677 not n20563 ; n20563_not
g39678 not n21139 ; n21139_not
g39679 not n22174 ; n22174_not
g39680 not n18313 ; n18313_not
g39681 not n17242 ; n17242_not
g39682 not n19150 ; n19150_not
g39683 not n22471 ; n22471_not
g39684 not n19141 ; n19141_not
g39685 not n21337 ; n21337_not
g39686 not n15352 ; n15352_not
g39687 not n21166 ; n21166_not
g39688 not n17251 ; n17251_not
g39689 not n22561 ; n22561_not
g39690 not n15343 ; n15343_not
g39691 not n20716 ; n20716_not
g39692 not n19213 ; n19213_not
g39693 not n18133 ; n18133_not
g39694 not n16801 ; n16801_not
g39695 not n19222 ; n19222_not
g39696 not n22552 ; n22552_not
g39697 not n21157 ; n21157_not
g39698 not n22255 ; n22255_not
g39699 not n19204 ; n19204_not
g39700 not n21904 ; n21904_not
g39701 not n22246 ; n22246_not
g39702 not n22543 ; n22543_not
g39703 not n17260 ; n17260_not
g39704 not n21148 ; n21148_not
g39705 not n20707 ; n20707_not
g39706 not n19231 ; n19231_not
g39707 not n20572 ; n20572_not
g39708 not n21346 ; n21346_not
g39709 not n19240 ; n19240_not
g39710 not n22291 ; n22291_not
g39711 not n18160 ; n18160_not
g39712 not n17314 ; n17314_not
g39713 not n20365 ; n20365_not
g39714 not n16342 ; n16342_not
g39715 not n15370 ; n15370_not
g39716 not n21418 ; n21418_not
g39717 not n20725 ; n20725_not
g39718 not n16135 ; n16135_not
g39719 not n22066 ; n22066_not
g39720 not n20086 ; n20086_not
g39721 not n22273 ; n22273_not
g39722 not n17305 ; n17305_not
g39723 not n20356 ; n20356_not
g39724 not n21850 ; n21850_not
g39725 not n20545 ; n20545_not
g39726 not n17332 ; n17332_not
g39727 not n20374 ; n20374_not
g39728 not n16522 ; n16522_not
g39729 not n16531 ; n16531_not
g39730 not n18520 ; n18520_not
g39731 not n16144 ; n16144_not
g39732 not n22804 ; n22804_not
g39733 not n21427 ; n21427_not
g39734 not n19402 ; n19402_not
g39735 not n15361 ; n15361_not
g39736 not n20842 ; n20842_not
g39737 not n17323 ; n17323_not
g39738 not n18331 ; n18331_not
g39739 not n21382 ; n21382_not
g39740 not n16360 ; n16360_not
g39741 not n18142 ; n18142_not
g39742 not n16504 ; n16504_not
g39743 not n22363 ; n22363_not
g39744 not n21364 ; n21364_not
g39745 not n16126 ; n16126_not
g39746 not n22057 ; n22057_not
g39747 not n22345 ; n22345_not
g39748 not n22570 ; n22570_not
g39749 not n18151 ; n18151_not
g39750 not n17620 ; n17620_not
g39751 not n16513 ; n16513_not
g39752 not n21409 ; n21409_not
g39753 not n22156 ; n22156_not
g39754 not n19321 ; n19321_not
g39755 not n20347 ; n20347_not
g39756 not n16900 ; n16900_not
g39757 not n20554 ; n20554_not
g39758 not n18403 ; n18403_not
g39759 not n19312 ; n19312_not
g39760 not n22606 ; n22606_not
g39761 not n16351 ; n16351_not
g39762 not n21391 ; n21391_not
g39763 not n18322 ; n18322_not
g39764 not n20338 ; n20338_not
g39765 not n17017 ; n17017_not
g39766 not n16018 ; n16018_not
g39767 not n18061 ; n18061_not
g39768 not n20950 ; n20950_not
g39769 not n15307 ; n15307_not
g39770 not n21229 ; n21229_not
g39771 not n20635 ; n20635_not
g39772 not n20095 ; n20095_not
g39773 not n17701 ; n17701_not
g39774 not n17161 ; n17161_not
g39775 not n16054 ; n16054_not
g39776 not n18052 ; n18052_not
g39777 not n22219 ; n22219_not
g39778 not n19015 ; n19015_not
g39779 not n27304 ; n27304_not
g39780 not n21265 ; n21265_not
g39781 not n17080 ; n17080_not
g39782 not n17170 ; n17170_not
g39783 not n17071 ; n17071_not
g39784 not n16063 ; n16063_not
g39785 not n15721 ; n15721_not
g39786 not n21274 ; n21274_not
g39787 not n16423 ; n16423_not
g39788 not n20617 ; n20617_not
g39789 not n20653 ; n20653_not
g39790 not n19033 ; n19033_not
g39791 not n18106 ; n18106_not
g39792 not n21283 ; n21283_not
g39793 not n18700 ; n18700_not
g39794 not n18601 ; n18601_not
g39795 not n20275 ; n20275_not
g39796 not n21247 ; n21247_not
g39797 not n20266 ; n20266_not
g39798 not n17125 ; n17125_not
g39799 not n20626 ; n20626_not
g39800 not n17134 ; n17134_not
g39801 not n18511 ; n18511_not
g39802 not n17116 ; n17116_not
g39803 not n15730 ; n15730_not
g39804 not n17107 ; n17107_not
g39805 not n23038 ; n23038_not
g39806 not n16036 ; n16036_not
g39807 not n18304 ; n18304_not
g39808 not n21238 ; n21238_not
g39809 not n16027 ; n16027_not
g39810 not n19006 ; n19006_not
g39811 not n17710 ; n17710_not
g39812 not n16405 ; n16405_not
g39813 not n20284 ; n20284_not
g39814 not n17143 ; n17143_not
g39815 not n17152 ; n17152_not
g39816 not n16045 ; n16045_not
g39817 not n16414 ; n16414_not
g39818 not n20257 ; n20257_not
g39819 not n22192 ; n22192_not
g39820 not n19114 ; n19114_not
g39821 not n21292 ; n21292_not
g39822 not n18016 ; n18016_not
g39823 not n15334 ; n15334_not
g39824 not n21940 ; n21940_not
g39825 not n20590 ; n20590_not
g39826 not n17215 ; n17215_not
g39827 not n22147 ; n22147_not
g39828 not n21184 ; n21184_not
g39829 not n16090 ; n16090_not
g39830 not n20680 ; n20680_not
g39831 not n18007 ; n18007_not
g39832 not n21706 ; n21706_not
g39833 not n20581 ; n20581_not
g39834 not n17224 ; n17224_not
g39835 not n21922 ; n21922_not
g39836 not n19132 ; n19132_not
g39837 not n15451 ; n15451_not
g39838 not n21913 ; n21913_not
g39839 not n22048 ; n22048_not
g39840 not n21319 ; n21319_not
g39841 not n22237 ; n22237_not
g39842 not n18124 ; n18124_not
g39843 not n22129 ; n22129_not
g39844 not n15253 ; n15253_not
g39845 not n17233 ; n17233_not
g39846 not n21049 ; n21049_not
g39847 not n17062 ; n17062_not
g39848 not n17521 ; n17521_not
g39849 not n18043 ; n18043_not
g39850 not n17053 ; n17053_not
g39851 not n19042 ; n19042_not
g39852 not n19051 ; n19051_not
g39853 not n17044 ; n17044_not
g39854 not n22525 ; n22525_not
g39855 not n18034 ; n18034_not
g39856 not n20608 ; n20608_not
g39857 not n16441 ; n16441_not
g39858 not n16009 ; n16009_not
g39859 not n16072 ; n16072_not
g39860 not n19060 ; n19060_not
g39861 not n22480 ; n22480_not
g39862 not n20662 ; n20662_not
g39863 not n15325 ; n15325_not
g39864 not n20671 ; n20671_not
g39865 not n22507 ; n22507_not
g39866 not n15712 ; n15712_not
g39867 not n18610 ; n18610_not
g39868 not n21193 ; n21193_not
g39869 not n17026 ; n17026_not
g39870 not n17206 ; n17206_not
g39871 not n22039 ; n22039_not
g39872 not n16081 ; n16081_not
g39873 not n17008 ; n17008_not
g39874 not n15604 ; n15604_not
g39875 not n18232 ; n18232_not
g39876 not n20464 ; n20464_not
g39877 not n21607 ; n21607_not
g39878 not n20806 ; n20806_not
g39879 not n22264 ; n22264_not
g39880 not n16234 ; n16234_not
g39881 not n21616 ; n21616_not
g39882 not n15505 ; n15505_not
g39883 not n20941 ; n20941_not
g39884 not n16603 ; n16603_not
g39885 not n20932 ; n20932_not
g39886 not n20158 ; n20158_not
g39887 not n20473 ; n20473_not
g39888 not n22390 ; n22390_not
g39889 not n15532 ; n15532_not
g39890 not n17503 ; n17503_not
g39891 not n22381 ; n22381_not
g39892 not n15523 ; n15523_not
g39893 not n16720 ; n16720_not
g39894 not n21625 ; n21625_not
g39895 not n16612 ; n16612_not
g39896 not n16243 ; n16243_not
g39897 not n15514 ; n15514_not
g39898 not n22426 ; n22426_not
g39899 not n15802 ; n15802_not
g39900 not n21535 ; n21535_not
g39901 not n18223 ; n18223_not
g39902 not n22831 ; n22831_not
g39903 not n17431 ; n17431_not
g39904 not n21724 ; n21724_not
g39905 not n21760 ; n21760_not
g39906 not n21544 ; n21544_not
g39907 not n15613 ; n15613_not
g39908 not n21553 ; n21553_not
g39909 not n21562 ; n21562_not
g39910 not n20176 ; n20176_not
g39911 not n16225 ; n16225_not
g39912 not n22354 ; n22354_not
g39913 not n17440 ; n17440_not
g39914 not n21751 ; n21751_not
g39915 not n16216 ; n16216_not
g39916 not n21472 ; n21472_not
g39917 not n22813 ; n22813_not
g39918 not n21571 ; n21571_not
g39919 not n21580 ; n21580_not
g39920 not n22822 ; n22822_not
g39921 not n17800 ; n17800_not
g39922 not n21661 ; n21661_not
g39923 not n22408 ; n22408_not
g39924 not n20491 ; n20491_not
g39925 not n22660 ; n22660_not
g39926 not n22723 ; n22723_not
g39927 not n17530 ; n17530_not
g39928 not n20860 ; n20860_not
g39929 not n21733 ; n21733_not
g39930 not n20851 ; n20851_not
g39931 not n22093 ; n22093_not
g39932 not n15811 ; n15811_not
g39933 not n20509 ; n20509_not
g39934 not n20833 ; n20833_not
g39935 not n17413 ; n17413_not
g39936 not n16630 ; n16630_not
g39937 not n21490 ; n21490_not
g39938 not n22417 ; n22417_not
g39939 not n22705 ; n22705_not
g39940 not n20518 ; n20518_not
g39941 not n20527 ; n20527_not
g39942 not n21715 ; n21715_not
g39943 not n20824 ; n20824_not
g39944 not n16261 ; n16261_not
g39945 not n22714 ; n22714_not
g39946 not n20059 ; n20059_not
g39947 not n16252 ; n16252_not
g39948 not n15091 ; n15091_not
g39949 not n20815 ; n20815_not
g39950 not n15550 ; n15550_not
g39951 not n22741 ; n22741_not
g39952 not n22750 ; n22750_not
g39953 not n15541 ; n15541_not
g39954 not n21643 ; n21643_not
g39955 not n20914 ; n20914_not
g39956 not n16702 ; n16702_not
g39957 not n21742 ; n21742_not
g39958 not n21634 ; n21634_not
g39959 not n20905 ; n20905_not
g39960 not n21670 ; n21670_not
g39961 not n18250 ; n18250_not
g39962 not n21652 ; n21652_not
g39963 not n20167 ; n20167_not
g39964 not n17512 ; n17512_not
g39965 not n18241 ; n18241_not
g39966 not n15208 ; n15208_not
g39967 not n18070 ; n18070_not
g39968 not n21058 ; n21058_not
g39969 not n20194 ; n20194_not
g39970 not n20392 ; n20392_not
g39971 not n22615 ; n22615_not
g39972 not n20077 ; n20077_not
g39973 not n22624 ; n22624_not
g39974 not n20734 ; n20734_not
g39975 not n21823 ; n21823_not
g39976 not n20743 ; n20743_not
g39977 not n19600 ; n19600_not
g39978 not n16333 ; n16333_not
g39979 not n19510 ; n19510_not
g39980 not n15910 ; n15910_not
g39981 not n22327 ; n22327_not
g39982 not n20068 ; n20068_not
g39983 not n22075 ; n22075_not
g39984 not n20185 ; n20185_not
g39985 not n21463 ; n21463_not
g39986 not n16171 ; n16171_not
g39987 not n15415 ; n15415_not
g39988 not n22318 ; n22318_not
g39989 not n21832 ; n21832_not
g39990 not n17341 ; n17341_not
g39991 not n19411 ; n19411_not
g39992 not n21841 ; n21841_not
g39993 not n22921 ; n22921_not
g39994 not n17350 ; n17350_not
g39995 not n21085 ; n21085_not
g39996 not n16153 ; n16153_not
g39997 not n22165 ; n22165_not
g39998 not n22444 ; n22444_not
g39999 not n22309 ; n22309_not
g40000 not n22462 ; n22462_not
g40001 not n18502 ; n18502_not
g40002 not n21067 ; n21067_not
g40003 not n20383 ; n20383_not
g40004 not n21076 ; n21076_not
g40005 not n16540 ; n16540_not
g40006 not n15406 ; n15406_not
g40007 not n21454 ; n21454_not
g40008 not n21445 ; n21445_not
g40009 not n21517 ; n21517_not
g40010 not n20536 ; n20536_not
g40011 not n17422 ; n17422_not
g40012 not n20437 ; n20437_not
g40013 not n20761 ; n20761_not
g40014 not n16315 ; n16315_not
g40015 not n15622 ; n15622_not
g40016 not n15280 ; n15280_not
g40017 not n16810 ; n16810_not
g40018 not n20329 ; n20329_not
g40019 not n18430 ; n18430_not
g40020 not n22138 ; n22138_not
g40021 not n22840 ; n22840_not
g40022 not n22642 ; n22642_not
g40023 not n20149 ; n20149_not
g40024 not n18412 ; n18412_not
g40025 not n21526 ; n21526_not
g40026 not n20446 ; n20446_not
g40027 not n20770 ; n20770_not
g40028 not n15460 ; n15460_not
g40029 not n18214 ; n18214_not
g40030 not n15640 ; n15640_not
g40031 not n17404 ; n17404_not
g40032 not n22336 ; n22336_not
g40033 not n16180 ; n16180_not
g40034 not n16306 ; n16306_not
g40035 not n15901 ; n15901_not
g40036 not n22435 ; n22435_not
g40037 not n21481 ; n21481_not
g40038 not n20428 ; n20428_not
g40039 not n22633 ; n22633_not
g40040 not n15433 ; n15433_not
g40041 not n18205 ; n18205_not
g40042 not n17602 ; n17602_not
g40043 not n15631 ; n15631_not
g40044 not n22903 ; n22903_not
g40045 not n16324 ; n16324_not
g40046 not n20419 ; n20419_not
g40047 not n21805 ; n21805_not
g40048 not n15424 ; n15424_not
g40049 not n21508 ; n21508_not
g40050 not n20752 ; n20752_not
g40051 not n26008 ; n26008_not
g40052 not n11590 ; n11590_not
g40053 not n25144 ; n25144_not
g40054 not n14614 ; n14614_not
g40055 not n23371 ; n23371_not
g40056 not n26125 ; n26125_not
g40057 not n14605 ; n14605_not
g40058 not n11608 ; n11608_not
g40059 not n25153 ; n25153_not
g40060 not n23605 ; n23605_not
g40061 not n14191 ; n14191_not
g40062 not n24253 ; n24253_not
g40063 not n11617 ; n11617_not
g40064 not n11626 ; n11626_not
g40065 not n25162 ; n25162_not
g40066 not n11248 ; n11248_not
g40067 not n11635 ; n11635_not
g40068 not n13804 ; n13804_not
g40069 not n14182 ; n14182_not
g40070 not n13741 ; n13741_not
g40071 not n11653 ; n11653_not
g40072 not n25171 ; n25171_not
g40073 not n12760 ; n12760_not
g40074 not n11509 ; n11509_not
g40075 not n11518 ; n11518_not
g40076 not n23560 ; n23560_not
g40077 not n25117 ; n25117_not
g40078 not n26170 ; n26170_not
g40079 not n26161 ; n26161_not
g40080 not n24280 ; n24280_not
g40081 not n11185 ; n11185_not
g40082 not n11527 ; n11527_not
g40083 not n11536 ; n11536_not
g40084 not n11545 ; n11545_not
g40085 not n12805 ; n12805_not
g40086 not n24271 ; n24271_not
g40087 not n14632 ; n14632_not
g40088 not n11554 ; n11554_not
g40089 not n26143 ; n26143_not
g40090 not n25126 ; n25126_not
g40091 not n14623 ; n14623_not
g40092 not n24073 ; n24073_not
g40093 not n11572 ; n11572_not
g40094 not n11563 ; n11563_not
g40095 not n25135 ; n25135_not
g40096 not n26134 ; n26134_not
g40097 not n11581 ; n11581_not
g40098 not n12715 ; n12715_not
g40099 not n14551 ; n14551_not
g40100 not n23461 ; n23461_not
g40101 not n11743 ; n11743_not
g40102 not n24226 ; n24226_not
g40103 not n26080 ; n26080_not
g40104 not n12706 ; n12706_not
g40105 not n13840 ; n13840_not
g40106 not n26071 ; n26071_not
g40107 not n25216 ; n25216_not
g40108 not n11752 ; n11752_not
g40109 not n12391 ; n12391_not
g40110 not n26062 ; n26062_not
g40111 not n11761 ; n11761_not
g40112 not n14542 ; n14542_not
g40113 not n26053 ; n26053_not
g40114 not n26044 ; n26044_not
g40115 not n25054 ; n25054_not
g40116 not n14533 ; n14533_not
g40117 not n12634 ; n12634_not
g40118 not n25225 ; n25225_not
g40119 not n24028 ; n24028_not
g40120 not n26116 ; n26116_not
g40121 not n25180 ; n25180_not
g40122 not n11671 ; n11671_not
g40123 not n11482 ; n11482_not
g40124 not n26107 ; n26107_not
g40125 not n23623 ; n23623_not
g40126 not n12751 ; n12751_not
g40127 not n13705 ; n13705_not
g40128 not n14164 ; n14164_not
g40129 not n23515 ; n23515_not
g40130 not n12733 ; n12733_not
g40131 not n23641 ; n23641_not
g40132 not n25207 ; n25207_not
g40133 not n11707 ; n11707_not
g40134 not n13822 ; n13822_not
g40135 not n11716 ; n11716_not
g40136 not n11725 ; n11725_not
g40137 not n24235 ; n24235_not
g40138 not n11329 ; n11329_not
g40139 not n14560 ; n14560_not
g40140 not n11734 ; n11734_not
g40141 not n13831 ; n13831_not
g40142 not n10843 ; n10843_not
g40143 not n23443 ; n23443_not
g40144 not n23452 ; n23452_not
g40145 not n24334 ; n24334_not
g40146 not n26242 ; n26242_not
g40147 not n13723 ; n13723_not
g40148 not n12931 ; n12931_not
g40149 not n13732 ; n13732_not
g40150 not n11158 ; n11158_not
g40151 not n12922 ; n12922_not
g40152 not n11266 ; n11266_not
g40153 not n26233 ; n26233_not
g40154 not n11275 ; n11275_not
g40155 not n14740 ; n14740_not
g40156 not n11284 ; n11284_not
g40157 not n12913 ; n12913_not
g40158 not n26224 ; n26224_not
g40159 not n11293 ; n11293_not
g40160 not n11338 ; n11338_not
g40161 not n25009 ; n25009_not
g40162 not n26260 ; n26260_not
g40163 not n23407 ; n23407_not
g40164 not n25018 ; n25018_not
g40165 not n23416 ; n23416_not
g40166 not n10717 ; n10717_not
g40167 not n11068 ; n11068_not
g40168 not n11086 ; n11086_not
g40169 not n23218 ; n23218_not
g40170 not n13714 ; n13714_not
g40171 not n23425 ; n23425_not
g40172 not n10933 ; n10933_not
g40173 not n23434 ; n23434_not
g40174 not n10852 ; n10852_not
g40175 not n12940 ; n12940_not
g40176 not n23182 ; n23182_not
g40177 not n11149 ; n11149_not
g40178 not n12562 ; n12562_not
g40179 not n11167 ; n11167_not
g40180 not n14731 ; n14731_not
g40181 not n23506 ; n23506_not
g40182 not n25090 ; n25090_not
g40183 not n26206 ; n26206_not
g40184 not n11419 ; n11419_not
g40185 not n11437 ; n11437_not
g40186 not n12850 ; n12850_not
g40187 not n11446 ; n11446_not
g40188 not n11383 ; n11383_not
g40189 not n11464 ; n11464_not
g40190 not n25108 ; n25108_not
g40191 not n11473 ; n11473_not
g40192 not n23524 ; n23524_not
g40193 not n12832 ; n12832_not
g40194 not n24307 ; n24307_not
g40195 not n23533 ; n23533_not
g40196 not n11491 ; n11491_not
g40197 not n12841 ; n12841_not
g40198 not n14650 ; n14650_not
g40199 not n23542 ; n23542_not
g40200 not n23551 ; n23551_not
g40201 not n12823 ; n12823_not
g40202 not n25036 ; n25036_not
g40203 not n14290 ; n14290_not
g40204 not n11347 ; n11347_not
g40205 not n11356 ; n11356_not
g40206 not n12616 ; n12616_not
g40207 not n11365 ; n11365_not
g40208 not n25063 ; n25063_not
g40209 not n24325 ; n24325_not
g40210 not n13750 ; n13750_not
g40211 not n11095 ; n11095_not
g40212 not n14713 ; n14713_not
g40213 not n25072 ; n25072_not
g40214 not n14704 ; n14704_not
g40215 not n25081 ; n25081_not
g40216 not n11392 ; n11392_not
g40217 not n26152 ; n26152_not
g40218 not n24316 ; n24316_not
g40219 not n12094 ; n12094_not
g40220 not n25522 ; n25522_not
g40221 not n12490 ; n12490_not
g40222 not n25351 ; n25351_not
g40223 not n12139 ; n12139_not
g40224 not n25513 ; n25513_not
g40225 not n14056 ; n14056_not
g40226 not n12148 ; n12148_not
g40227 not n12481 ; n12481_not
g40228 not n25360 ; n25360_not
g40229 not n12166 ; n12166_not
g40230 not n24082 ; n24082_not
g40231 not n14236 ; n14236_not
g40232 not n12175 ; n12175_not
g40233 not n14065 ; n14065_not
g40234 not n12184 ; n12184_not
g40235 not n11815 ; n11815_not
g40236 not n14254 ; n14254_not
g40237 not n25504 ; n25504_not
g40238 not n12193 ; n12193_not
g40239 not n14245 ; n14245_not
g40240 not n25540 ; n25540_not
g40241 not n14344 ; n14344_not
g40242 not n23902 ; n23902_not
g40243 not n14335 ; n14335_not
g40244 not n25531 ; n25531_not
g40245 not n12049 ; n12049_not
g40246 not n14029 ; n14029_not
g40247 not n12058 ; n12058_not
g40248 not n14326 ; n14326_not
g40249 not n12067 ; n12067_not
g40250 not n14317 ; n14317_not
g40251 not n12076 ; n12076_not
g40252 not n14308 ; n14308_not
g40253 not n14038 ; n14038_not
g40254 not n23911 ; n23911_not
g40255 not n23920 ; n23920_not
g40256 not n12085 ; n12085_not
g40257 not n14047 ; n14047_not
g40258 not n12409 ; n12409_not
g40259 not n24037 ; n24037_not
g40260 not n14083 ; n14083_not
g40261 not n12337 ; n12337_not
g40262 not n12328 ; n12328_not
g40263 not n11941 ; n11941_not
g40264 not n12346 ; n12346_not
g40265 not n14173 ; n14173_not
g40266 not n24064 ; n24064_not
g40267 not n25414 ; n25414_not
g40268 not n25432 ; n25432_not
g40269 not n24055 ; n24055_not
g40270 not n12355 ; n12355_not
g40271 not n14155 ; n14155_not
g40272 not n12382 ; n12382_not
g40273 not n14119 ; n14119_not
g40274 not n12364 ; n12364_not
g40275 not n14146 ; n14146_not
g40276 not n25423 ; n25423_not
g40277 not n14137 ; n14137_not
g40278 not n12373 ; n12373_not
g40279 not n14128 ; n14128_not
g40280 not n14074 ; n14074_not
g40281 not n12472 ; n12472_not
g40282 not n12238 ; n12238_not
g40283 not n23812 ; n23812_not
g40284 not n12463 ; n12463_not
g40285 not n12247 ; n12247_not
g40286 not n25342 ; n25342_not
g40287 not n12256 ; n12256_not
g40288 not n14209 ; n14209_not
g40289 not n12265 ; n12265_not
g40290 not n12274 ; n12274_not
g40291 not n12454 ; n12454_not
g40292 not n24019 ; n24019_not
g40293 not n12436 ; n12436_not
g40294 not n12292 ; n12292_not
g40295 not n25441 ; n25441_not
g40296 not n12418 ; n12418_not
g40297 not n12319 ; n12319_not
g40298 not n11842 ; n11842_not
g40299 not n25900 ; n25900_not
g40300 not n23740 ; n23740_not
g40301 not n11851 ; n11851_not
g40302 not n24163 ; n24163_not
g40303 not n25810 ; n25810_not
g40304 not n11860 ; n11860_not
g40305 not n25252 ; n25252_not
g40306 not n24172 ; n24172_not
g40307 not n13912 ; n13912_not
g40308 not n23632 ; n23632_not
g40309 not n12643 ; n12643_not
g40310 not n14470 ; n14470_not
g40311 not n14461 ; n14461_not
g40312 not n13921 ; n13921_not
g40313 not n25261 ; n25261_not
g40314 not n14218 ; n14218_not
g40315 not n27241 ; n27241_not
g40316 not n25270 ; n25270_not
g40317 not n23803 ; n23803_not
g40318 not n25234 ; n25234_not
g40319 not n23704 ; n23704_not
g40320 not n11770 ; n11770_not
g40321 not n14515 ; n14515_not
g40322 not n24208 ; n24208_not
g40323 not n26026 ; n26026_not
g40324 not n14506 ; n14506_not
g40325 not n11455 ; n11455_not
g40326 not n11806 ; n11806_not
g40327 not n23713 ; n23713_not
g40328 not n24190 ; n24190_not
g40329 not n23722 ; n23722_not
g40330 not n11824 ; n11824_not
g40331 not n12661 ; n12661_not
g40332 not n25243 ; n25243_not
g40333 not n24181 ; n24181_not
g40334 not n23731 ; n23731_not
g40335 not n25324 ; n25324_not
g40336 not n12544 ; n12544_not
g40337 not n24118 ; n24118_not
g40338 not n23821 ; n23821_not
g40339 not n24109 ; n24109_not
g40340 not n25630 ; n25630_not
g40341 not n13570 ; n13570_not
g40342 not n12535 ; n12535_not
g40343 not n24091 ; n24091_not
g40344 not n25621 ; n25621_not
g40345 not n14380 ; n14380_not
g40346 not n25612 ; n25612_not
g40347 not n14371 ; n14371_not
g40348 not n12526 ; n12526_not
g40349 not n25603 ; n25603_not
g40350 not n12517 ; n12517_not
g40351 not n12508 ; n12508_not
g40352 not n14362 ; n14362_not
g40353 not n14443 ; n14443_not
g40354 not n25801 ; n25801_not
g40355 not n24154 ; n24154_not
g40356 not n12580 ; n12580_not
g40357 not n11905 ; n11905_not
g40358 not n25306 ; n25306_not
g40359 not n12571 ; n12571_not
g40360 not n14425 ; n14425_not
g40361 not n25315 ; n25315_not
g40362 not n12229 ; n12229_not
g40363 not n25720 ; n25720_not
g40364 not n25711 ; n25711_not
g40365 not n14416 ; n14416_not
g40366 not n14407 ; n14407_not
g40367 not n24136 ; n24136_not
g40368 not n24127 ; n24127_not
g40369 not n25702 ; n25702_not
g40370 not n11950 ; n11950_not
g40371 not n27043 ; n27043_not
g40372 not n13606 ; n13606_not
g40373 not n10582 ; n10582_not
g40374 not n23128 ; n23128_not
g40375 not n10591 ; n10591_not
g40376 not n15136 ; n15136_not
g40377 not n23245 ; n23245_not
g40378 not n13390 ; n13390_not
g40379 not n15145 ; n15145_not
g40380 not n13615 ; n13615_not
g40381 not n26800 ; n26800_not
g40382 not n26710 ; n26710_not
g40383 not n15154 ; n15154_not
g40384 not n10618 ; n10618_not
g40385 not n13255 ; n13255_not
g40386 not n10636 ; n10636_not
g40387 not n14920 ; n14920_not
g40388 not n10537 ; n10537_not
g40389 not n15118 ; n15118_not
g40390 not n10555 ; n10555_not
g40391 not n13147 ; n13147_not
g40392 not n13273 ; n13273_not
g40393 not n24604 ; n24604_not
g40394 not n10564 ; n10564_not
g40395 not n13381 ; n13381_not
g40396 not n23227 ; n23227_not
g40397 not n15127 ; n15127_not
g40398 not n10573 ; n10573_not
g40399 not n10087 ; n10087_not
g40400 not n10069 ; n10069_not
g40401 not n24424 ; n24424_not
g40402 not n10672 ; n10672_not
g40403 not n10690 ; n10690_not
g40404 not n13192 ; n13192_not
g40405 not n15172 ; n15172_not
g40406 not n26422 ; n26422_not
g40407 not n14902 ; n14902_not
g40408 not n26620 ; n26620_not
g40409 not n13183 ; n13183_not
g40410 not n13426 ; n13426_not
g40411 not n26611 ; n26611_not
g40412 not n24550 ; n24550_not
g40413 not n10663 ; n10663_not
g40414 not n13246 ; n13246_not
g40415 not n10726 ; n10726_not
g40416 not n24712 ; n24712_not
g40417 not n24415 ; n24415_not
g40418 not n10735 ; n10735_not
g40419 not n27232 ; n27232_not
g40420 not n10645 ; n10645_not
g40421 not n10654 ; n10654_not
g40422 not n13408 ; n13408_not
g40423 not n23119 ; n23119_not
g40424 not n15163 ; n15163_not
g40425 not n13552 ; n13552_not
g40426 not n23263 ; n23263_not
g40427 not n12904 ; n12904_not
g40428 not n13624 ; n13624_not
g40429 not n13237 ; n13237_not
g40430 not n27250 ; n27250_not
g40431 not n23272 ; n23272_not
g40432 not n13219 ; n13219_not
g40433 not n26701 ; n26701_not
g40434 not n10681 ; n10681_not
g40435 not n24703 ; n24703_not
g40436 not n14830 ; n14830_not
g40437 not n23155 ; n23155_not
g40438 not n13354 ; n13354_not
g40439 not n15037 ; n15037_not
g40440 not n13309 ; n13309_not
g40441 not n24433 ; n24433_not
g40442 not n24460 ; n24460_not
g40443 not n27025 ; n27025_not
g40444 not n10339 ; n10339_not
g40445 not n15082 ; n15082_not
g40446 not n10348 ; n10348_not
g40447 not n15019 ; n15019_not
g40448 not n24631 ; n24631_not
g40449 not n10249 ; n10249_not
g40450 not n24451 ; n24451_not
g40451 not n10276 ; n10276_not
g40452 not n10195 ; n10195_not
g40453 not n10357 ; n10357_not
g40454 not n24613 ; n24613_not
g40455 not n10366 ; n10366_not
g40456 not n10186 ; n10186_not
g40457 not n23146 ; n23146_not
g40458 not n13336 ; n13336_not
g40459 not n15073 ; n15073_not
g40460 not n13345 ; n13345_not
g40461 not n13327 ; n13327_not
g40462 not n10285 ; n10285_not
g40463 not n15064 ; n15064_not
g40464 not n27034 ; n27034_not
g40465 not n23137 ; n23137_not
g40466 not n10267 ; n10267_not
g40467 not n24622 ; n24622_not
g40468 not n10258 ; n10258_not
g40469 not n10294 ; n10294_not
g40470 not n15046 ; n15046_not
g40471 not n13318 ; n13318_not
g40472 not n10456 ; n10456_not
g40473 not n23191 ; n23191_not
g40474 not n10078 ; n10078_not
g40475 not n13282 ; n13282_not
g40476 not n10465 ; n10465_not
g40477 not n27007 ; n27007_not
g40478 not n10483 ; n10483_not
g40479 not n10492 ; n10492_not
g40480 not n13372 ; n13372_not
g40481 not n23209 ; n23209_not
g40482 not n10168 ; n10168_not
g40483 not n10519 ; n10519_not
g40484 not n15109 ; n15109_not
g40485 not n10528 ; n10528_not
g40486 not n10375 ; n10375_not
g40487 not n13291 ; n13291_not
g40488 not n23056 ; n23056_not
g40489 not n10177 ; n10177_not
g40490 not n23164 ; n23164_not
g40491 not n23173 ; n23173_not
g40492 not n10429 ; n10429_not
g40493 not n10393 ; n10393_not
g40494 not n27016 ; n27016_not
g40495 not n10438 ; n10438_not
g40496 not n10447 ; n10447_not
g40497 not n13651 ; n13651_not
g40498 not n15244 ; n15244_not
g40499 not n10834 ; n10834_not
g40500 not n13075 ; n13075_not
g40501 not n27313 ; n27313_not
g40502 not n23344 ; n23344_not
g40503 not n13264 ; n13264_not
g40504 not n13462 ; n13462_not
g40505 not n24406 ; n24406_not
g40506 not n26503 ; n26503_not
g40507 not n10942 ; n10942_not
g40508 not n10780 ; n10780_not
g40509 not n24820 ; n24820_not
g40510 not n10807 ; n10807_not
g40511 not n23326 ; n23326_not
g40512 not n24532 ; n24532_not
g40513 not n15055 ; n15055_not
g40514 not n23335 ; n23335_not
g40515 not n15235 ; n15235_not
g40516 not n24514 ; n24514_not
g40517 not n24541 ; n24541_not
g40518 not n10960 ; n10960_not
g40519 not n10816 ; n10816_not
g40520 not n24505 ; n24505_not
g40521 not n24901 ; n24901_not
g40522 not n10825 ; n10825_not
g40523 not n26341 ; n26341_not
g40524 not n13039 ; n13039_not
g40525 not n27115 ; n27115_not
g40526 not n24811 ; n24811_not
g40527 not n26413 ; n26413_not
g40528 not n13480 ; n13480_not
g40529 not n26404 ; n26404_not
g40530 not n15271 ; n15271_not
g40531 not n23362 ; n23362_not
g40532 not n13435 ; n13435_not
g40533 not n23074 ; n23074_not
g40534 not n27142 ; n27142_not
g40535 not n23065 ; n23065_not
g40536 not n15262 ; n15262_not
g40537 not n24370 ; n24370_not
g40538 not n24523 ; n24523_not
g40539 not n10861 ; n10861_not
g40540 not n13066 ; n13066_not
g40541 not n26440 ; n26440_not
g40542 not n13057 ; n13057_not
g40543 not n13471 ; n13471_not
g40544 not n10753 ; n10753_not
g40545 not n14812 ; n14812_not
g40546 not n13048 ; n13048_not
g40547 not n13660 ; n13660_not
g40548 not n26350 ; n26350_not
g40549 not n13174 ; n13174_not
g40550 not n27070 ; n27070_not
g40551 not n10762 ; n10762_not
g40552 not n13516 ; n13516_not
g40553 not n27124 ; n27124_not
g40554 not n24910 ; n24910_not
g40555 not n27223 ; n27223_not
g40556 not n27106 ; n27106_not
g40557 not n13165 ; n13165_not
g40558 not n23083 ; n23083_not
g40559 not n10771 ; n10771_not
g40560 not n24244 ; n24244_not
g40561 not n13507 ; n13507_not
g40562 not n15190 ; n15190_not
g40563 not n24361 ; n24361_not
g40564 not n23281 ; n23281_not
g40565 not n23047 ; n23047_not
g40566 not n10744 ; n10744_not
g40567 not n13543 ; n13543_not
g40568 not n26602 ; n26602_not
g40569 not n27061 ; n27061_not
g40570 not n23317 ; n23317_not
g40571 not n13633 ; n13633_not
g40572 not n13444 ; n13444_not
g40573 not n24730 ; n24730_not
g40574 not n26314 ; n26314_not
g40575 not n15217 ; n15217_not
g40576 not n27205 ; n27205_not
g40577 not n15226 ; n15226_not
g40578 not n13642 ; n13642_not
g40579 not n13534 ; n13534_not
g40580 not n23380 ; n23380_not
g40581 not n24217 ; n24217_not
g40582 not n26512 ; n26512_not
g40583 not n26323 ; n26323_not
g40584 not n13093 ; n13093_not
g40585 not n13138 ; n13138_not
g40586 not n13129 ; n13129_not
g40587 not n26530 ; n26530_not
g40588 not n12536 ; n12536_not
g40589 not n13490 ; n13490_not
g40590 not n13337 ; n13337_not
g40591 not n16730 ; n16730_not
g40592 not n25325 ; n25325_not
g40593 not n13481 ; n13481_not
g40594 not n17306 ; n17306_not
g40595 not n16721 ; n16721_not
g40596 not n12554 ; n12554_not
g40597 not n13364 ; n13364_not
g40598 not n12392 ; n12392_not
g40599 not n13355 ; n13355_not
g40600 not n25316 ; n25316_not
g40601 not n25415 ; n25415_not
g40602 not n17315 ; n17315_not
g40603 not n12266 ; n12266_not
g40604 not n12563 ; n12563_not
g40605 not n21185 ; n21185_not
g40606 not n21626 ; n21626_not
g40607 not n21725 ; n21725_not
g40608 not n13346 ; n13346_not
g40609 not n24614 ; n24614_not
g40610 not n21743 ; n21743_not
g40611 not n17225 ; n17225_not
g40612 not n24524 ; n24524_not
g40613 not n13382 ; n13382_not
g40614 not n25343 ; n25343_not
g40615 not n21644 ; n21644_not
g40616 not n21653 ; n21653_not
g40617 not n24560 ; n24560_not
g40618 not n24542 ; n24542_not
g40619 not n21662 ; n21662_not
g40620 not n25370 ; n25370_not
g40621 not n21671 ; n21671_not
g40622 not n13409 ; n13409_not
g40623 not n16640 ; n16640_not
g40624 not n17243 ; n17243_not
g40625 not n25361 ; n25361_not
g40626 not n20870 ; n20870_not
g40627 not n21446 ; n21446_not
g40628 not n13418 ; n13418_not
g40629 not n12482 ; n12482_not
g40630 not n17270 ; n17270_not
g40631 not n25352 ; n25352_not
g40632 not n24551 ; n24551_not
g40633 not n21680 ; n21680_not
g40634 not n13445 ; n13445_not
g40635 not n12491 ; n12491_not
g40636 not n12473 ; n12473_not
g40637 not n21149 ; n21149_not
g40638 not n24425 ; n24425_not
g40639 not n21635 ; n21635_not
g40640 not n12518 ; n12518_not
g40641 not n13094 ; n13094_not
g40642 not n12527 ; n12527_not
g40643 not n21086 ; n21086_not
g40644 not n16622 ; n16622_not
g40645 not n21167 ; n21167_not
g40646 not n13373 ; n13373_not
g40647 not n21176 ; n21176_not
g40648 not n17234 ; n17234_not
g40649 not n16712 ; n16712_not
g40650 not n16613 ; n16613_not
g40651 not n25406 ; n25406_not
g40652 not n24227 ; n24227_not
g40653 not n25163 ; n25163_not
g40654 not n12455 ; n12455_not
g40655 not n12437 ; n12437_not
g40656 not n13463 ; n13463_not
g40657 not n16631 ; n16631_not
g40658 not n16703 ; n16703_not
g40659 not n21158 ; n21158_not
g40660 not n24605 ; n24605_not
g40661 not n12509 ; n12509_not
g40662 not n24533 ; n24533_not
g40663 not n16343 ; n16343_not
g40664 not n12428 ; n12428_not
g40665 not n12419 ; n12419_not
g40666 not n13166 ; n13166_not
g40667 not n12824 ; n12824_not
g40668 not n21293 ; n21293_not
g40669 not n13148 ; n13148_not
g40670 not n17036 ; n17036_not
g40671 not n12833 ; n12833_not
g40672 not n25109 ; n25109_not
g40673 not n21455 ; n21455_not
g40674 not n17027 ; n17027_not
g40675 not n12842 ; n12842_not
g40676 not n24731 ; n24731_not
g40677 not n17018 ; n17018_not
g40678 not n12851 ; n12851_not
g40679 not n25091 ; n25091_not
g40680 not n13085 ; n13085_not
g40681 not n12860 ; n12860_not
g40682 not n17009 ; n17009_not
g40683 not n13076 ; n13076_not
g40684 not n25145 ; n25145_not
g40685 not n17072 ; n17072_not
g40686 not n25136 ; n25136_not
g40687 not n24704 ; n24704_not
g40688 not n13184 ; n13184_not
g40689 not n21275 ; n21275_not
g40690 not n25127 ; n25127_not
g40691 not n17063 ; n17063_not
g40692 not n12671 ; n12671_not
g40693 not n21284 ; n21284_not
g40694 not n21491 ; n21491_not
g40695 not n17054 ; n17054_not
g40696 not n12806 ; n12806_not
g40697 not n21194 ; n21194_not
g40698 not n25118 ; n25118_not
g40699 not n24713 ; n24713_not
g40700 not n17045 ; n17045_not
g40701 not n12815 ; n12815_not
g40702 not n21482 ; n21482_not
g40703 not n21329 ; n21329_not
g40704 not n12932 ; n12932_not
g40705 not n12590 ; n12590_not
g40706 not n21392 ; n21392_not
g40707 not n21374 ; n21374_not
g40708 not n24821 ; n24821_not
g40709 not n16910 ; n16910_not
g40710 not n21338 ; n21338_not
g40711 not n25028 ; n25028_not
g40712 not n21383 ; n21383_not
g40713 not n24902 ; n24902_not
g40714 not n12941 ; n12941_not
g40715 not n21068 ; n21068_not
g40716 not n25019 ; n25019_not
g40717 not n12950 ; n12950_not
g40718 not n24911 ; n24911_not
g40719 not n24830 ; n24830_not
g40720 not n21356 ; n21356_not
g40721 not n25082 ; n25082_not
g40722 not n21428 ; n21428_not
g40723 not n25073 ; n25073_not
g40724 not n13067 ; n13067_not
g40725 not n25055 ; n25055_not
g40726 not n13058 ; n13058_not
g40727 not n12905 ; n12905_not
g40728 not n25037 ; n25037_not
g40729 not n13049 ; n13049_not
g40730 not n24803 ; n24803_not
g40731 not n12914 ; n12914_not
g40732 not n24812 ; n24812_not
g40733 not n16901 ; n16901_not
g40734 not n12923 ; n12923_not
g40735 not n24623 ; n24623_not
g40736 not n12653 ; n12653_not
g40737 not n25253 ; n25253_not
g40738 not n13292 ; n13292_not
g40739 not n17162 ; n17162_not
g40740 not n21590 ; n21590_not
g40741 not n25244 ; n25244_not
g40742 not n16604 ; n16604_not
g40743 not n12662 ; n12662_not
g40744 not n25226 ; n25226_not
g40745 not n24632 ; n24632_not
g40746 not n21581 ; n21581_not
g40747 not n17153 ; n17153_not
g40748 not n21572 ; n21572_not
g40749 not n13283 ; n13283_not
g40750 not n21239 ; n21239_not
g40751 not n25235 ; n25235_not
g40752 not n21563 ; n21563_not
g40753 not n12680 ; n12680_not
g40754 not n17207 ; n17207_not
g40755 not n12572 ; n12572_not
g40756 not n13328 ; n13328_not
g40757 not n25307 ; n25307_not
g40758 not n12581 ; n12581_not
g40759 not n25280 ; n25280_not
g40760 not n13319 ; n13319_not
g40761 not n21608 ; n21608_not
g40762 not n25271 ; n25271_not
g40763 not n12617 ; n12617_not
g40764 not n25262 ; n25262_not
g40765 not n17180 ; n17180_not
g40766 not n12635 ; n12635_not
g40767 not n12644 ; n12644_not
g40768 not n17171 ; n17171_not
g40769 not n16802 ; n16802_not
g40770 not n25208 ; n25208_not
g40771 not n24470 ; n24470_not
g40772 not n21527 ; n21527_not
g40773 not n12734 ; n12734_not
g40774 not n25190 ; n25190_not
g40775 not n13256 ; n13256_not
g40776 not n25181 ; n25181_not
g40777 not n21248 ; n21248_not
g40778 not n13238 ; n13238_not
g40779 not n17090 ; n17090_not
g40780 not n21257 ; n21257_not
g40781 not n16811 ; n16811_not
g40782 not n21518 ; n21518_not
g40783 not n13229 ; n13229_not
g40784 not n16235 ; n16235_not
g40785 not n12770 ; n12770_not
g40786 not n25154 ; n25154_not
g40787 not n21266 ; n21266_not
g40788 not n16820 ; n16820_not
g40789 not n13193 ; n13193_not
g40790 not n17135 ; n17135_not
g40791 not n21554 ; n21554_not
g40792 not n25217 ; n25217_not
g40793 not n17126 ; n17126_not
g40794 not n21473 ; n21473_not
g40795 not n21545 ; n21545_not
g40796 not n24641 ; n24641_not
g40797 not n16280 ; n16280_not
g40798 not n13274 ; n13274_not
g40799 not n12707 ; n12707_not
g40800 not n17108 ; n17108_not
g40801 not n17117 ; n17117_not
g40802 not n21536 ; n21536_not
g40803 not n12716 ; n12716_not
g40804 not n12725 ; n12725_not
g40805 not n24650 ; n24650_not
g40806 not n13265 ; n13265_not
g40807 not n13247 ; n13247_not
g40808 not n10817 ; n10817_not
g40809 not n10808 ; n10808_not
g40810 not n18206 ; n18206_not
g40811 not n10448 ; n10448_not
g40812 not n10790 ; n10790_not
g40813 not n18215 ; n18215_not
g40814 not n26513 ; n26513_not
g40815 not n20177 ; n20177_not
g40816 not n26522 ; n26522_not
g40817 not n10781 ; n10781_not
g40818 not n18224 ; n18224_not
g40819 not n26531 ; n26531_not
g40820 not n18233 ; n18233_not
g40821 not n26450 ; n26450_not
g40822 not n26423 ; n26423_not
g40823 not n18152 ; n18152_not
g40824 not n18071 ; n18071_not
g40825 not n10862 ; n10862_not
g40826 not n18170 ; n18170_not
g40827 not n10853 ; n10853_not
g40828 not n10844 ; n10844_not
g40829 not n20195 ; n20195_not
g40830 not n26504 ; n26504_not
g40831 not n10835 ; n10835_not
g40832 not n20186 ; n20186_not
g40833 not n26621 ; n26621_not
g40834 not n10691 ; n10691_not
g40835 not n26603 ; n26603_not
g40836 not n26540 ; n26540_not
g40837 not n10682 ; n10682_not
g40838 not n26702 ; n26702_not
g40839 not n18035 ; n18035_not
g40840 not n10673 ; n10673_not
g40841 not n26711 ; n26711_not
g40842 not n10664 ; n10664_not
g40843 not n26720 ; n26720_not
g40844 not n10655 ; n10655_not
g40845 not n18305 ; n18305_not
g40846 not n10619 ; n10619_not
g40847 not n18242 ; n18242_not
g40848 not n10763 ; n10763_not
g40849 not n20168 ; n20168_not
g40850 not n18251 ; n18251_not
g40851 not n20159 ; n20159_not
g40852 not n18260 ; n18260_not
g40853 not n10736 ; n10736_not
g40854 not n10727 ; n10727_not
g40855 not n10718 ; n10718_not
g40856 not n26612 ; n26612_not
g40857 not n10709 ; n10709_not
g40858 not n11177 ; n11177_not
g40859 not n11168 ; n11168_not
g40860 not n18017 ; n18017_not
g40861 not n26243 ; n26243_not
g40862 not n18026 ; n18026_not
g40863 not n26252 ; n26252_not
g40864 not n11096 ; n11096_not
g40865 not n11087 ; n11087_not
g40866 not n11078 ; n11078_not
g40867 not n11069 ; n11069_not
g40868 not n18044 ; n18044_not
g40869 not n18053 ; n18053_not
g40870 not n26135 ; n26135_not
g40871 not n26261 ; n26261_not
g40872 not n20348 ; n20348_not
g40873 not n17630 ; n17630_not
g40874 not n11348 ; n11348_not
g40875 not n11339 ; n11339_not
g40876 not n20339 ; n20339_not
g40877 not n11294 ; n11294_not
g40878 not n11285 ; n11285_not
g40879 not n11267 ; n11267_not
g40880 not n11249 ; n11249_not
g40881 not n11159 ; n11159_not
g40882 not n10826 ; n10826_not
g40883 not n26234 ; n26234_not
g40884 not n26225 ; n26225_not
g40885 not n11195 ; n11195_not
g40886 not n11186 ; n11186_not
g40887 not n26342 ; n26342_not
g40888 not n10934 ; n10934_not
g40889 not n26351 ; n26351_not
g40890 not n26360 ; n26360_not
g40891 not n10916 ; n10916_not
g40892 not n10754 ; n10754_not
g40893 not n18125 ; n18125_not
g40894 not n10907 ; n10907_not
g40895 not n26405 ; n26405_not
g40896 not n18143 ; n18143_not
g40897 not n10880 ; n10880_not
g40898 not n26414 ; n26414_not
g40899 not n18062 ; n18062_not
g40900 not n20285 ; n20285_not
g40901 not n26270 ; n26270_not
g40902 not n26216 ; n26216_not
g40903 not n20276 ; n20276_not
g40904 not n26306 ; n26306_not
g40905 not n18080 ; n18080_not
g40906 not n20267 ; n20267_not
g40907 not n26315 ; n26315_not
g40908 not n20258 ; n20258_not
g40909 not n10961 ; n10961_not
g40910 not n26324 ; n26324_not
g40911 not n10952 ; n10952_not
g40912 not n18107 ; n18107_not
g40913 not n27260 ; n27260_not
g40914 not n19223 ; n19223_not
g40915 not n27251 ; n27251_not
g40916 not n19214 ; n19214_not
g40917 not n19205 ; n19205_not
g40918 not n27242 ; n27242_not
g40919 not n19160 ; n19160_not
g40920 not n19151 ; n19151_not
g40921 not n27233 ; n27233_not
g40922 not n19070 ; n19070_not
g40923 not n27224 ; n27224_not
g40924 not n10178 ; n10178_not
g40925 not n18521 ; n18521_not
g40926 not n18512 ; n18512_not
g40927 not n10079 ; n10079_not
g40928 not n10169 ; n10169_not
g40929 not n18530 ; n18530_not
g40930 not n19340 ; n19340_not
g40931 not n27044 ; n27044_not
g40932 not n19322 ; n19322_not
g40933 not n10097 ; n10097_not
g40934 not n10088 ; n10088_not
g40935 not n19304 ; n19304_not
g40936 not n27008 ; n27008_not
g40937 not n19034 ; n19034_not
g40938 not n19241 ; n19241_not
g40939 not n19232 ; n19232_not
g40940 not n27161 ; n27161_not
g40941 not n19016 ; n19016_not
g40942 not n27125 ; n27125_not
g40943 not n27143 ; n27143_not
g40944 not n19007 ; n19007_not
g40945 not n27107 ; n27107_not
g40946 not n27071 ; n27071_not
g40947 not n27116 ; n27116_not
g40948 not n18332 ; n18332_not
g40949 not n27134 ; n27134_not
g40950 not n18800 ; n18800_not
g40951 not n18431 ; n18431_not
g40952 not n18701 ; n18701_not
g40953 not n27062 ; n27062_not
g40954 not n18602 ; n18602_not
g40955 not n19115 ; n19115_not
g40956 not n27206 ; n27206_not
g40957 not n27152 ; n27152_not
g40958 not n19106 ; n19106_not
g40959 not n18620 ; n18620_not
g40960 not n27080 ; n27080_not
g40961 not n18611 ; n18611_not
g40962 not n19061 ; n19061_not
g40963 not n19052 ; n19052_not
g40964 not n19043 ; n19043_not
g40965 not n10196 ; n10196_not
g40966 not n10538 ; n10538_not
g40967 not n10529 ; n10529_not
g40968 not n10187 ; n10187_not
g40969 not n10466 ; n10466_not
g40970 not n10367 ; n10367_not
g40971 not n10457 ; n10457_not
g40972 not n10439 ; n10439_not
g40973 not n27017 ; n27017_not
g40974 not n10394 ; n10394_not
g40975 not n20096 ; n20096_not
g40976 not n26810 ; n26810_not
g40977 not n10592 ; n10592_not
g40978 not n20087 ; n20087_not
g40979 not n10583 ; n10583_not
g40980 not n26900 ; n26900_not
g40981 not n18341 ; n18341_not
g40982 not n20078 ; n20078_not
g40983 not n10574 ; n10574_not
g40984 not n20069 ; n20069_not
g40985 not n18350 ; n18350_not
g40986 not n10556 ; n10556_not
g40987 not n10547 ; n10547_not
g40988 not n10277 ; n10277_not
g40989 not n19601 ; n19601_not
g40990 not n10268 ; n10268_not
g40991 not n19403 ; n19403_not
g40992 not n19520 ; n19520_not
g40993 not n19511 ; n19511_not
g40994 not n10259 ; n10259_not
g40995 not n19502 ; n19502_not
g40996 not n19430 ; n19430_not
g40997 not n18503 ; n18503_not
g40998 not n19412 ; n19412_not
g40999 not n18404 ; n18404_not
g41000 not n10376 ; n10376_not
g41001 not n18413 ; n18413_not
g41002 not n27026 ; n27026_not
g41003 not n18422 ; n18422_not
g41004 not n10358 ; n10358_not
g41005 not n10349 ; n10349_not
g41006 not n10286 ; n10286_not
g41007 not n10295 ; n10295_not
g41008 not n18440 ; n18440_not
g41009 not n19700 ; n19700_not
g41010 not n17531 ; n17531_not
g41011 not n17540 ; n17540_not
g41012 not n20861 ; n20861_not
g41013 not n20852 ; n20852_not
g41014 not n25703 ; n25703_not
g41015 not n20843 ; n20843_not
g41016 not n11942 ; n11942_not
g41017 not n20834 ; n20834_not
g41018 not n25712 ; n25712_not
g41019 not n25721 ; n25721_not
g41020 not n25730 ; n25730_not
g41021 not n11924 ; n11924_not
g41022 not n20816 ; n20816_not
g41023 not n25604 ; n25604_not
g41024 not n17504 ; n17504_not
g41025 not n20915 ; n20915_not
g41026 not n25613 ; n25613_not
g41027 not n20681 ; n20681_not
g41028 not n17144 ; n17144_not
g41029 not n25622 ; n25622_not
g41030 not n17513 ; n17513_not
g41031 not n17360 ; n17360_not
g41032 not n25514 ; n25514_not
g41033 not n20906 ; n20906_not
g41034 not n11960 ; n11960_not
g41035 not n25640 ; n25640_not
g41036 not n25820 ; n25820_not
g41037 not n20744 ; n20744_not
g41038 not n20663 ; n20663_not
g41039 not n17612 ; n17612_not
g41040 not n20735 ; n20735_not
g41041 not n11870 ; n11870_not
g41042 not n20726 ; n20726_not
g41043 not n25901 ; n25901_not
g41044 not n25910 ; n25910_not
g41045 not n25631 ; n25631_not
g41046 not n20807 ; n20807_not
g41047 not n11915 ; n11915_not
g41048 not n11906 ; n11906_not
g41049 not n20780 ; n20780_not
g41050 not n20771 ; n20771_not
g41051 not n25802 ; n25802_not
g41052 not n20762 ; n20762_not
g41053 not n20627 ; n20627_not
g41054 not n25811 ; n25811_not
g41055 not n20753 ; n20753_not
g41056 not n17603 ; n17603_not
g41057 not n21077 ; n21077_not
g41058 not n25442 ; n25442_not
g41059 not n12293 ; n12293_not
g41060 not n11618 ; n11618_not
g41061 not n25460 ; n25460_not
g41062 not n21059 ; n21059_not
g41063 not n12275 ; n12275_not
g41064 not n12248 ; n12248_not
g41065 not n12239 ; n12239_not
g41066 not n12149 ; n12149_not
g41067 not n12185 ; n12185_not
g41068 not n12167 ; n12167_not
g41069 not n25505 ; n25505_not
g41070 not n12374 ; n12374_not
g41071 not n12365 ; n12365_not
g41072 not n25424 ; n25424_not
g41073 not n12356 ; n12356_not
g41074 not n17333 ; n17333_not
g41075 not n21095 ; n21095_not
g41076 not n25433 ; n25433_not
g41077 not n17342 ; n17342_not
g41078 not n12347 ; n12347_not
g41079 not n12338 ; n12338_not
g41080 not n12329 ; n12329_not
g41081 not n12077 ; n12077_not
g41082 not n17450 ; n17450_not
g41083 not n12059 ; n12059_not
g41084 not n11852 ; n11852_not
g41085 not n25532 ; n25532_not
g41086 not n25541 ; n25541_not
g41087 not n20960 ; n20960_not
g41088 not n25550 ; n25550_not
g41089 not n20951 ; n20951_not
g41090 not n20933 ; n20933_not
g41091 not n25451 ; n25451_not
g41092 not n12176 ; n12176_not
g41093 not n17414 ; n17414_not
g41094 not n12158 ; n12158_not
g41095 not n17423 ; n17423_not
g41096 not n11816 ; n11816_not
g41097 not n17432 ; n17432_not
g41098 not n25523 ; n25523_not
g41099 not n12095 ; n12095_not
g41100 not n17441 ; n17441_not
g41101 not n12086 ; n12086_not
g41102 not n20474 ; n20474_not
g41103 not n20465 ; n20465_not
g41104 not n26153 ; n26153_not
g41105 not n11546 ; n11546_not
g41106 not n20456 ; n20456_not
g41107 not n11537 ; n11537_not
g41108 not n20447 ; n20447_not
g41109 not n11528 ; n11528_not
g41110 not n26162 ; n26162_not
g41111 not n26171 ; n26171_not
g41112 not n11519 ; n11519_not
g41113 not n17900 ; n17900_not
g41114 not n20438 ; n20438_not
g41115 not n11636 ; n11636_not
g41116 not n11627 ; n11627_not
g41117 not n11483 ; n11483_not
g41118 not n11609 ; n11609_not
g41119 not n20519 ; n20519_not
g41120 not n26126 ; n26126_not
g41121 not n11582 ; n11582_not
g41122 not n11591 ; n11591_not
g41123 not n20492 ; n20492_not
g41124 not n20483 ; n20483_not
g41125 not n11573 ; n11573_not
g41126 not n11564 ; n11564_not
g41127 not n20384 ; n20384_not
g41128 not n20393 ; n20393_not
g41129 not n11393 ; n11393_not
g41130 not n11384 ; n11384_not
g41131 not n20375 ; n20375_not
g41132 not n11375 ; n11375_not
g41133 not n20366 ; n20366_not
g41134 not n17621 ; n17621_not
g41135 not n20357 ; n20357_not
g41136 not n11357 ; n11357_not
g41137 not n20429 ; n20429_not
g41138 not n11492 ; n11492_not
g41139 not n26180 ; n26180_not
g41140 not n11474 ; n11474_not
g41141 not n11465 ; n11465_not
g41142 not n11456 ; n11456_not
g41143 not n11438 ; n11438_not
g41144 not n26207 ; n26207_not
g41145 not n26036 ; n26036_not
g41146 not n17702 ; n17702_not
g41147 not n20636 ; n20636_not
g41148 not n11780 ; n11780_not
g41149 not n26045 ; n26045_not
g41150 not n17711 ; n17711_not
g41151 not n11771 ; n11771_not
g41152 not n17720 ; n17720_not
g41153 not n26063 ; n26063_not
g41154 not n11762 ; n11762_not
g41155 not n20618 ; n20618_not
g41156 not n11753 ; n11753_not
g41157 not n20717 ; n20717_not
g41158 not n11843 ; n11843_not
g41159 not n11744 ; n11744_not
g41160 not n20708 ; n20708_not
g41161 not n11834 ; n11834_not
g41162 not n26009 ; n26009_not
g41163 not n20690 ; n20690_not
g41164 not n11825 ; n11825_not
g41165 not n20672 ; n20672_not
g41166 not n11807 ; n11807_not
g41167 not n26018 ; n26018_not
g41168 not n26027 ; n26027_not
g41169 not n20654 ; n20654_not
g41170 not n26090 ; n26090_not
g41171 not n11690 ; n11690_not
g41172 not n20546 ; n20546_not
g41173 not n26054 ; n26054_not
g41174 not n26108 ; n26108_not
g41175 not n20528 ; n20528_not
g41176 not n11672 ; n11672_not
g41177 not n17801 ; n17801_not
g41178 not n26117 ; n26117_not
g41179 not n11654 ; n11654_not
g41180 not n17810 ; n17810_not
g41181 not n11645 ; n11645_not
g41182 not n26072 ; n26072_not
g41183 not n20609 ; n20609_not
g41184 not n26081 ; n26081_not
g41185 not n20591 ; n20591_not
g41186 not n11735 ; n11735_not
g41187 not n20582 ; n20582_not
g41188 not n11726 ; n11726_not
g41189 not n20564 ; n20564_not
g41190 not n11708 ; n11708_not
g41191 not n20555 ; n20555_not
g41192 not n16046 ; n16046_not
g41193 not n23921 ; n23921_not
g41194 not n14291 ; n14291_not
g41195 not n16037 ; n16037_not
g41196 not n23912 ; n23912_not
g41197 not n14309 ; n14309_not
g41198 not n16028 ; n16028_not
g41199 not n16019 ; n16019_not
g41200 not n14327 ; n14327_not
g41201 not n23903 ; n23903_not
g41202 not n14345 ; n14345_not
g41203 not n14336 ; n14336_not
g41204 not n14354 ; n14354_not
g41205 not n14363 ; n14363_not
g41206 not n15614 ; n15614_not
g41207 not n23840 ; n23840_not
g41208 not n22229 ; n22229_not
g41209 not n14381 ; n14381_not
g41210 not n23831 ; n23831_not
g41211 not n22238 ; n22238_not
g41212 not n23732 ; n23732_not
g41213 not n23822 ; n23822_not
g41214 not n16109 ; n16109_not
g41215 not n14165 ; n14165_not
g41216 not n24038 ; n24038_not
g41217 not n14174 ; n14174_not
g41218 not n24029 ; n24029_not
g41219 not n15722 ; n15722_not
g41220 not n14183 ; n14183_not
g41221 not n16091 ; n16091_not
g41222 not n14192 ; n14192_not
g41223 not n14129 ; n14129_not
g41224 not n22193 ; n22193_not
g41225 not n16082 ; n16082_not
g41226 not n14057 ; n14057_not
g41227 not n13940 ; n13940_not
g41228 not n16073 ; n16073_not
g41229 not n14237 ; n14237_not
g41230 not n14246 ; n14246_not
g41231 not n14255 ; n14255_not
g41232 not n14264 ; n14264_not
g41233 not n14273 ; n14273_not
g41234 not n16055 ; n16055_not
g41235 not n23930 ; n23930_not
g41236 not n23741 ; n23741_not
g41237 not n14480 ; n14480_not
g41238 not n22337 ; n22337_not
g41239 not n15902 ; n15902_not
g41240 not n23723 ; n23723_not
g41241 not n22058 ; n22058_not
g41242 not n14507 ; n14507_not
g41243 not n22346 ; n22346_not
g41244 not n14516 ; n14516_not
g41245 not n23705 ; n23705_not
g41246 not n22355 ; n22355_not
g41247 not n22265 ; n22265_not
g41248 not n15542 ; n15542_not
g41249 not n15605 ; n15605_not
g41250 not n22364 ; n22364_not
g41251 not n14543 ; n14543_not
g41252 not n22382 ; n22382_not
g41253 not n23660 ; n23660_not
g41254 not n14147 ; n14147_not
g41255 not n14552 ; n14552_not
g41256 not n14561 ; n14561_not
g41257 not n22409 ; n22409_not
g41258 not n23642 ; n23642_not
g41259 not n14390 ; n14390_not
g41260 not n23813 ; n23813_not
g41261 not n22247 ; n22247_not
g41262 not n22256 ; n22256_not
g41263 not n14219 ; n14219_not
g41264 not n14417 ; n14417_not
g41265 not n14426 ; n14426_not
g41266 not n22274 ; n22274_not
g41267 not n14435 ; n14435_not
g41268 not n23804 ; n23804_not
g41269 not n22292 ; n22292_not
g41270 not n14444 ; n14444_not
g41271 not n23750 ; n23750_not
g41272 not n22319 ; n22319_not
g41273 not n15920 ; n15920_not
g41274 not n23633 ; n23633_not
g41275 not n15911 ; n15911_not
g41276 not n22328 ; n22328_not
g41277 not n16334 ; n16334_not
g41278 not n22076 ; n22076_not
g41279 not n16325 ; n16325_not
g41280 not n24272 ; n24272_not
g41281 not n16316 ; n16316_not
g41282 not n24263 ; n24263_not
g41283 not n24254 ; n24254_not
g41284 not n16307 ; n16307_not
g41285 not n24245 ; n24245_not
g41286 not n13805 ; n13805_not
g41287 not n22085 ; n22085_not
g41288 not n13823 ; n13823_not
g41289 not n22094 ; n22094_not
g41290 not n13841 ; n13841_not
g41291 not n16262 ; n16262_not
g41292 not n24209 ; n24209_not
g41293 not n24191 ; n24191_not
g41294 not n13706 ; n13706_not
g41295 not n24344 ; n24344_not
g41296 not n13715 ; n13715_not
g41297 not n24335 ; n24335_not
g41298 not n13724 ; n13724_not
g41299 not n24119 ; n24119_not
g41300 not n13733 ; n13733_not
g41301 not n16370 ; n16370_not
g41302 not n24326 ; n24326_not
g41303 not n13742 ; n13742_not
g41304 not n16361 ; n16361_not
g41305 not n13751 ; n13751_not
g41306 not n24317 ; n24317_not
g41307 not n16352 ; n16352_not
g41308 not n13760 ; n13760_not
g41309 not n22067 ; n22067_not
g41310 not n24308 ; n24308_not
g41311 not n24281 ; n24281_not
g41312 not n24290 ; n24290_not
g41313 not n22148 ; n22148_not
g41314 not n16181 ; n16181_not
g41315 not n24074 ; n24074_not
g41316 not n24083 ; n24083_not
g41317 not n16172 ; n16172_not
g41318 not n14039 ; n14039_not
g41319 not n22157 ; n22157_not
g41320 not n14048 ; n14048_not
g41321 not n13634 ; n13634_not
g41322 not n16154 ; n16154_not
g41323 not n14066 ; n14066_not
g41324 not n22166 ; n22166_not
g41325 not n14075 ; n14075_not
g41326 not n16136 ; n16136_not
g41327 not n14084 ; n14084_not
g41328 not n14093 ; n14093_not
g41329 not n24056 ; n24056_not
g41330 not n16127 ; n16127_not
g41331 not n13832 ; n13832_not
g41332 not n16118 ; n16118_not
g41333 not n16253 ; n16253_not
g41334 not n24182 ; n24182_not
g41335 not n16244 ; n16244_not
g41336 not n13904 ; n13904_not
g41337 not n24173 ; n24173_not
g41338 not n13913 ; n13913_not
g41339 not n24164 ; n24164_not
g41340 not n13922 ; n13922_not
g41341 not n13931 ; n13931_not
g41342 not n16226 ; n16226_not
g41343 not n24155 ; n24155_not
g41344 not n24146 ; n24146_not
g41345 not n16217 ; n16217_not
g41346 not n15830 ; n15830_not
g41347 not n13526 ; n13526_not
g41348 not n24137 ; n24137_not
g41349 not n24128 ; n24128_not
g41350 not n24092 ; n24092_not
g41351 not n16190 ; n16190_not
g41352 not n24065 ; n24065_not
g41353 not n23219 ; n23219_not
g41354 not n22841 ; n22841_not
g41355 not n22850 ; n22850_not
g41356 not n15461 ; n15461_not
g41357 not n15452 ; n15452_not
g41358 not n23192 ; n23192_not
g41359 not n22715 ; n22715_not
g41360 not n15443 ; n15443_not
g41361 not n23183 ; n23183_not
g41362 not n15434 ; n15434_not
g41363 not n23174 ; n23174_not
g41364 not n27314 ; n27314_not
g41365 not n15425 ; n15425_not
g41366 not n22904 ; n22904_not
g41367 not n14912 ; n14912_not
g41368 not n22670 ; n22670_not
g41369 not n15416 ; n15416_not
g41370 not n23156 ; n23156_not
g41371 not n15038 ; n15038_not
g41372 not n15029 ; n15029_not
g41373 not n15407 ; n15407_not
g41374 not n15056 ; n15056_not
g41375 not n22742 ; n22742_not
g41376 not n14408 ; n14408_not
g41377 not n23282 ; n23282_not
g41378 not n23066 ; n23066_not
g41379 not n22760 ; n22760_not
g41380 not n22751 ; n22751_not
g41381 not n15533 ; n15533_not
g41382 not n14903 ; n14903_not
g41383 not n23273 ; n23273_not
g41384 not n15524 ; n15524_not
g41385 not n23264 ; n23264_not
g41386 not n15515 ; n15515_not
g41387 not n23255 ; n23255_not
g41388 not n14921 ; n14921_not
g41389 not n23246 ; n23246_not
g41390 not n23165 ; n23165_not
g41391 not n22814 ; n22814_not
g41392 not n23237 ; n23237_not
g41393 not n23228 ; n23228_not
g41394 not n15470 ; n15470_not
g41395 not n22832 ; n22832_not
g41396 not n15344 ; n15344_not
g41397 not n15173 ; n15173_not
g41398 not n15191 ; n15191_not
g41399 not n23093 ; n23093_not
g41400 not n23084 ; n23084_not
g41401 not n15209 ; n15209_not
g41402 not n15326 ; n15326_not
g41403 not n15218 ; n15218_not
g41404 not n15227 ; n15227_not
g41405 not n15236 ; n15236_not
g41406 not n15317 ; n15317_not
g41407 not n23075 ; n23075_not
g41408 not n15254 ; n15254_not
g41409 not n15308 ; n15308_not
g41410 not n15263 ; n15263_not
g41411 not n15272 ; n15272_not
g41412 not n23057 ; n23057_not
g41413 not n14651 ; n14651_not
g41414 not n23039 ; n23039_not
g41415 not n15281 ; n15281_not
g41416 not n23048 ; n23048_not
g41417 not n15290 ; n15290_not
g41418 not n15065 ; n15065_not
g41419 not n15074 ; n15074_not
g41420 not n22922 ; n22922_not
g41421 not n22940 ; n22940_not
g41422 not n15083 ; n15083_not
g41423 not n15380 ; n15380_not
g41424 not n22913 ; n22913_not
g41425 not n23138 ; n23138_not
g41426 not n15371 ; n15371_not
g41427 not n15119 ; n15119_not
g41428 not n23129 ; n23129_not
g41429 not n15362 ; n15362_not
g41430 not n15128 ; n15128_not
g41431 not n15137 ; n15137_not
g41432 not n15146 ; n15146_not
g41433 not n15353 ; n15353_not
g41434 not n15155 ; n15155_not
g41435 not n15164 ; n15164_not
g41436 not n23543 ; n23543_not
g41437 not n23534 ; n23534_not
g41438 not n22508 ; n22508_not
g41439 not n14660 ; n14660_not
g41440 not n15740 ; n15740_not
g41441 not n23525 ; n23525_not
g41442 not n22517 ; n22517_not
g41443 not n15731 ; n15731_not
g41444 not n23516 ; n23516_not
g41445 not n22526 ; n22526_not
g41446 not n23480 ; n23480_not
g41447 not n15713 ; n15713_not
g41448 not n14705 ; n14705_not
g41449 not n14714 ; n14714_not
g41450 not n23471 ; n23471_not
g41451 not n22544 ; n22544_not
g41452 not n14732 ; n14732_not
g41453 not n23435 ; n23435_not
g41454 not n23624 ; n23624_not
g41455 not n22418 ; n22418_not
g41456 not n14570 ; n14570_not
g41457 not n15812 ; n15812_not
g41458 not n23615 ; n23615_not
g41459 not n22427 ; n22427_not
g41460 not n23552 ; n23552_not
g41461 not n15803 ; n15803_not
g41462 not n22184 ; n22184_not
g41463 not n23606 ; n23606_not
g41464 not n22436 ; n22436_not
g41465 not n14606 ; n14606_not
g41466 not n14615 ; n14615_not
g41467 not n22445 ; n22445_not
g41468 not n14624 ; n14624_not
g41469 not n23561 ; n23561_not
g41470 not n22472 ; n22472_not
g41471 not n14633 ; n14633_not
g41472 not n22481 ; n22481_not
g41473 not n22490 ; n22490_not
g41474 not n15506 ; n15506_not
g41475 not n23363 ; n23363_not
g41476 not n14831 ; n14831_not
g41477 not n22661 ; n22661_not
g41478 not n23345 ; n23345_not
g41479 not n14840 ; n14840_not
g41480 not n22706 ; n22706_not
g41481 not n23336 ; n23336_not
g41482 not n23327 ; n23327_not
g41483 not n23318 ; n23318_not
g41484 not n22724 ; n22724_not
g41485 not n15560 ; n15560_not
g41486 not n23291 ; n23291_not
g41487 not n15551 ; n15551_not
g41488 not n22562 ; n22562_not
g41489 not n22580 ; n22580_not
g41490 not n27305 ; n27305_not
g41491 not n22463 ; n22463_not
g41492 not n23453 ; n23453_not
g41493 not n14750 ; n14750_not
g41494 not n23444 ; n23444_not
g41495 not n22616 ; n22616_not
g41496 not n15650 ; n15650_not
g41497 not n23417 ; n23417_not
g41498 not n22625 ; n22625_not
g41499 not n23408 ; n23408_not
g41500 not n15641 ; n15641_not
g41501 not n15632 ; n15632_not
g41502 not n23381 ; n23381_not
g41503 not n22634 ; n22634_not
g41504 not n14804 ; n14804_not
g41505 not n15623 ; n15623_not
g41506 not n23372 ; n23372_not
g41507 not n14813 ; n14813_not
g41508 not n22643 ; n22643_not
g41509 not n24407 ; n24407_not
g41510 not n13472 ; n13472_not
g41511 not n24218 ; n24218_not
g41512 not n24434 ; n24434_not
g41513 not n24371 ; n24371_not
g41514 not n21851 ; n21851_not
g41515 not n21806 ; n21806_not
g41516 not n21914 ; n21914_not
g41517 not n21860 ; n21860_not
g41518 not n21905 ; n21905_not
g41519 not n16433 ; n16433_not
g41520 not n21815 ; n21815_not
g41521 not n16415 ; n16415_not
g41522 not n13643 ; n13643_not
g41523 not n13616 ; n13616_not
g41524 not n13625 ; n13625_not
g41525 not n16406 ; n16406_not
g41526 not n13535 ; n13535_not
g41527 not n13661 ; n13661_not
g41528 not n16523 ; n16523_not
g41529 not n16541 ; n16541_not
g41530 not n13508 ; n13508_not
g41531 not n24362 ; n24362_not
g41532 not n21770 ; n21770_not
g41533 not n13571 ; n13571_not
g41534 not n13436 ; n13436_not
g41535 not n21752 ; n21752_not
g41536 not n16532 ; n16532_not
g41537 not n13553 ; n13553_not
g41538 not n13607 ; n13607_not
g41539 not n21932 ; n21932_not
g41540 not n24461 ; n24461_not
g41541 not n24506 ; n24506_not
g41542 not n24353 ; n24353_not
g41543 not n21707 ; n21707_not
g41544 not n24416 ; n24416_not
g41545 not n21842 ; n21842_not
g41546 not n24380 ; n24380_not
g41547 not n13517 ; n13517_not
g41548 not n16514 ; n16514_not
g41549 not n13670 ; n13670_not
g41550 not n21761 ; n21761_not
g41551 not n16460 ; n16460_not
g41552 not n21824 ; n21824_not
g41553 not n13544 ; n13544_not
g41554 not n21950 ; n21950_not
g41555 not n16424 ; n16424_not
g41556 not n13652 ; n13652_not
g41557 not n21941 ; n21941_not
g41558 not n16442 ; n16442_not
g41559 not n21833 ; n21833_not
g41560 not n11574 ; n11574_not
g41561 not n19710 ; n19710_not
g41562 not n20484 ; n20484_not
g41563 not n16506 ; n16506_not
g41564 not n11592 ; n11592_not
g41565 not n14616 ; n14616_not
g41566 not n11484 ; n11484_not
g41567 not n22455 ; n22455_not
g41568 not n19530 ; n19530_not
g41569 not n22446 ; n22446_not
g41570 not n20493 ; n20493_not
g41571 not n19800 ; n19800_not
g41572 not n24633 ; n24633_not
g41573 not n23580 ; n23580_not
g41574 not n11583 ; n11583_not
g41575 not n26136 ; n26136_not
g41576 not n16461 ; n16461_not
g41577 not n10287 ; n10287_not
g41578 not n11637 ; n11637_not
g41579 not n22185 ; n22185_not
g41580 not n17811 ; n17811_not
g41581 not n19341 ; n19341_not
g41582 not n11646 ; n11646_not
g41583 not n23616 ; n23616_not
g41584 not n21807 ; n21807_not
g41585 not n11655 ; n11655_not
g41586 not n26118 ; n26118_not
g41587 not n11664 ; n11664_not
g41588 not n14580 ; n14580_not
g41589 not n15813 ; n15813_not
g41590 not n17802 ; n17802_not
g41591 not n16173 ; n16173_not
g41592 not n20538 ; n20538_not
g41593 not n11673 ; n11673_not
g41594 not n19701 ; n19701_not
g41595 not n18450 ; n18450_not
g41596 not n15057 ; n15057_not
g41597 not n26127 ; n26127_not
g41598 not n21573 ; n21573_not
g41599 not n18108 ; n18108_not
g41600 not n22437 ; n22437_not
g41601 not n24435 ; n24435_not
g41602 not n15408 ; n15408_not
g41603 not n22194 ; n22194_not
g41604 not n21564 ; n21564_not
g41605 not n15435 ; n15435_not
g41606 not n11619 ; n11619_not
g41607 not n13590 ; n13590_not
g41608 not n11628 ; n11628_not
g41609 not n17820 ; n17820_not
g41610 not n15804 ; n15804_not
g41611 not n24273 ; n24273_not
g41612 not n22428 ; n22428_not
g41613 not n14661 ; n14661_not
g41614 not n11475 ; n11475_not
g41615 not n15327 ; n15327_not
g41616 not n26181 ; n26181_not
g41617 not n11367 ; n11367_not
g41618 not n13293 ; n13293_not
g41619 not n13581 ; n13581_not
g41620 not n26073 ; n26073_not
g41621 not n22905 ; n22905_not
g41622 not n22509 ; n22509_not
g41623 not n21591 ; n21591_not
g41624 not n17910 ; n17910_not
g41625 not n21861 ; n21861_not
g41626 not n23535 ; n23535_not
g41627 not n11493 ; n11493_not
g41628 not n16650 ; n16650_not
g41629 not n26172 ; n26172_not
g41630 not n17901 ; n17901_not
g41631 not n24453 ; n24453_not
g41632 not n15723 ; n15723_not
g41633 not n26208 ; n26208_not
g41634 not n26163 ; n26163_not
g41635 not n18414 ; n18414_not
g41636 not n15426 ; n15426_not
g41637 not n23517 ; n23517_not
g41638 not n13437 ; n13437_not
g41639 not n22518 ; n22518_not
g41640 not n11439 ; n11439_not
g41641 not n16641 ; n16641_not
g41642 not n18423 ; n18423_not
g41643 not n10359 ; n10359_not
g41644 not n11457 ; n11457_not
g41645 not n15732 ; n15732_not
g41646 not n26190 ; n26190_not
g41647 not n13284 ; n13284_not
g41648 not n16560 ; n16560_not
g41649 not n22473 ; n22473_not
g41650 not n11538 ; n11538_not
g41651 not n20457 ; n20457_not
g41652 not n13446 ; n13446_not
g41653 not n24444 ; n24444_not
g41654 not n22464 ; n22464_not
g41655 not n11547 ; n11547_not
g41656 not n23562 ; n23562_not
g41657 not n22356 ; n22356_not
g41658 not n20466 ; n20466_not
g41659 not n26154 ; n26154_not
g41660 not n11556 ; n11556_not
g41661 not n11565 ; n11565_not
g41662 not n23571 ; n23571_not
g41663 not n15039 ; n15039_not
g41664 not n20475 ; n20475_not
g41665 not n14625 ; n14625_not
g41666 not n20439 ; n20439_not
g41667 not n15750 ; n15750_not
g41668 not n23553 ; n23553_not
g41669 not n14643 ; n14643_not
g41670 not n21582 ; n21582_not
g41671 not n27027 ; n27027_not
g41672 not n22491 ; n22491_not
g41673 not n15390 ; n15390_not
g41674 not n17514 ; n17514_not
g41675 not n15417 ; n15417_not
g41676 not n22293 ; n22293_not
g41677 not n11529 ; n11529_not
g41678 not n23157 ; n23157_not
g41679 not n22482 ; n22482_not
g41680 not n20448 ; n20448_not
g41681 not n23328 ; n23328_not
g41682 not n18432 ; n18432_not
g41683 not n14634 ; n14634_not
g41684 not n10296 ; n10296_not
g41685 not n19422 ; n19422_not
g41686 not n14481 ; n14481_not
g41687 not n11835 ; n11835_not
g41688 not n24651 ; n24651_not
g41689 not n19413 ; n19413_not
g41690 not n20709 ; n20709_not
g41691 not n15903 ; n15903_not
g41692 not n11844 ; n11844_not
g41693 not n10188 ; n10188_not
g41694 not n16803 ; n16803_not
g41695 not n25911 ; n25911_not
g41696 not n13608 ; n13608_not
g41697 not n20718 ; n20718_not
g41698 not n23742 ; n23742_not
g41699 not n15381 ; n15381_not
g41700 not n16263 ; n16263_not
g41701 not n17640 ; n17640_not
g41702 not n13257 ; n13257_not
g41703 not n23733 ; n23733_not
g41704 not n18513 ; n18513_not
g41705 not n15084 ; n15084_not
g41706 not n14508 ; n14508_not
g41707 not n11466 ; n11466_not
g41708 not n10197 ; n10197_not
g41709 not n22347 ; n22347_not
g41710 not n23634 ; n23634_not
g41711 not n11808 ; n11808_not
g41712 not n22950 ; n22950_not
g41713 not n26019 ; n26019_not
g41714 not n23715 ; n23715_not
g41715 not n20673 ; n20673_not
g41716 not n14490 ; n14490_not
g41717 not n18504 ; n18504_not
g41718 not n20358 ; n20358_not
g41719 not n11817 ; n11817_not
g41720 not n19206 ; n19206_not
g41721 not n22338 ; n22338_not
g41722 not n20682 ; n20682_not
g41723 not n21906 ; n21906_not
g41724 not n23724 ; n23724_not
g41725 not n20691 ; n20691_not
g41726 not n11826 ; n11826_not
g41727 not n20664 ; n20664_not
g41728 not n22914 ; n22914_not
g41729 not n25830 ; n25830_not
g41730 not n25812 ; n25812_not
g41731 not n17613 ; n17613_not
g41732 not n24660 ; n24660_not
g41733 not n19404 ; n19404_not
g41734 not n14463 ; n14463_not
g41735 not n20745 ; n20745_not
g41736 not n25821 ; n25821_not
g41737 not n23760 ; n23760_not
g41738 not n21726 ; n21726_not
g41739 not n15372 ; n15372_not
g41740 not n17604 ; n17604_not
g41741 not n15930 ; n15930_not
g41742 not n23607 ; n23607_not
g41743 not n14454 ; n14454_not
g41744 not n14445 ; n14445_not
g41745 not n12861 ; n12861_not
g41746 not n20754 ; n20754_not
g41747 not n13239 ; n13239_not
g41748 not n13464 ; n13464_not
g41749 not n25920 ; n25920_not
g41750 not n17631 ; n17631_not
g41751 not n15912 ; n15912_not
g41752 not n17622 ; n17622_not
g41753 not n21915 ; n21915_not
g41754 not n13248 ; n13248_not
g41755 not n10179 ; n10179_not
g41756 not n25902 ; n25902_not
g41757 not n15921 ; n15921_not
g41758 not n22266 ; n22266_not
g41759 not n11871 ; n11871_not
g41760 not n23751 ; n23751_not
g41761 not n20736 ; n20736_not
g41762 not n13617 ; n13617_not
g41763 not n20727 ; n20727_not
g41764 not n18522 ; n18522_not
g41765 not n10269 ; n10269_not
g41766 not n15075 ; n15075_not
g41767 not n23643 ; n23643_not
g41768 not n20565 ; n20565_not
g41769 not n15840 ; n15840_not
g41770 not n14562 ; n14562_not
g41771 not n11727 ; n11727_not
g41772 not n26082 ; n26082_not
g41773 not n13266 ; n13266_not
g41774 not n17451 ; n17451_not
g41775 not n20583 ; n20583_not
g41776 not n23652 ; n23652_not
g41777 not n20592 ; n20592_not
g41778 not n19521 ; n19521_not
g41779 not n22383 ; n22383_not
g41780 not n11745 ; n11745_not
g41781 not n13275 ; n13275_not
g41782 not n19620 ; n19620_not
g41783 not n21870 ; n21870_not
g41784 not n15822 ; n15822_not
g41785 not n26109 ; n26109_not
g41786 not n24642 ; n24642_not
g41787 not n11682 ; n11682_not
g41788 not n22419 ; n22419_not
g41789 not n22923 ; n22923_not
g41790 not n14571 ; n14571_not
g41791 not n20547 ; n20547_not
g41792 not n24543 ; n24543_not
g41793 not n26055 ; n26055_not
g41794 not n11691 ; n11691_not
g41795 not n26091 ; n26091_not
g41796 not n19611 ; n19611_not
g41797 not n20556 ; n20556_not
g41798 not n21546 ; n21546_not
g41799 not n11709 ; n11709_not
g41800 not n22239 ; n22239_not
g41801 not n13455 ; n13455_not
g41802 not n17712 ; n17712_not
g41803 not n26046 ; n26046_not
g41804 not n23670 ; n23670_not
g41805 not n21537 ; n21537_not
g41806 not n20637 ; n20637_not
g41807 not n19440 ; n19440_not
g41808 not n17334 ; n17334_not
g41809 not n14526 ; n14526_not
g41810 not n17703 ; n17703_not
g41811 not n14517 ; n14517_not
g41812 not n11781 ; n11781_not
g41813 not n19431 ; n19431_not
g41814 not n26037 ; n26037_not
g41815 not n20646 ; n20646_not
g41816 not n27036 ; n27036_not
g41817 not n26028 ; n26028_not
g41818 not n11790 ; n11790_not
g41819 not n23706 ; n23706_not
g41820 not n20655 ; n20655_not
g41821 not n23661 ; n23661_not
g41822 not n19512 ; n19512_not
g41823 not n11754 ; n11754_not
g41824 not n19503 ; n19503_not
g41825 not n22374 ; n22374_not
g41826 not n20619 ; n20619_not
g41827 not n26064 ; n26064_not
g41828 not n14544 ; n14544_not
g41829 not n17730 ; n17730_not
g41830 not n21528 ; n21528_not
g41831 not n22365 ; n22365_not
g41832 not n15633 ; n15633_not
g41833 not n11763 ; n11763_not
g41834 not n17721 ; n17721_not
g41835 not n21708 ; n21708_not
g41836 not n22932 ; n22932_not
g41837 not n14535 ; n14535_not
g41838 not n11772 ; n11772_not
g41839 not n13527 ; n13527_not
g41840 not n27315 ; n27315_not
g41841 not n10845 ; n10845_not
g41842 not n10791 ; n10791_not
g41843 not n21834 ; n21834_not
g41844 not n26442 ; n26442_not
g41845 not n22815 ; n22815_not
g41846 not n26820 ; n26820_not
g41847 not n22671 ; n22671_not
g41848 not n26460 ; n26460_not
g41849 not n21672 ; n21672_not
g41850 not n13374 ; n13374_not
g41851 not n10854 ; n10854_not
g41852 not n18333 ; n18333_not
g41853 not n18171 ; n18171_not
g41854 not n26406 ; n26406_not
g41855 not n26451 ; n26451_not
g41856 not n23346 ; n23346_not
g41857 not n15480 ; n15480_not
g41858 not n23238 ; n23238_not
g41859 not n18342 ; n18342_not
g41860 not n10863 ; n10863_not
g41861 not n10575 ; n10575_not
g41862 not n18207 ; n18207_not
g41863 not n22635 ; n22635_not
g41864 not n23337 ; n23337_not
g41865 not n13563 ; n13563_not
g41866 not n10818 ; n10818_not
g41867 not n10809 ; n10809_not
g41868 not n22707 ; n22707_not
g41869 not n10827 ; n10827_not
g41870 not n20187 ; n20187_not
g41871 not n18018 ; n18018_not
g41872 not n10584 ; n10584_not
g41873 not n14850 ; n14850_not
g41874 not n10836 ; n10836_not
g41875 not n14841 ; n14841_not
g41876 not n26505 ; n26505_not
g41877 not n16704 ; n16704_not
g41878 not n15570 ; n15570_not
g41879 not n20196 ; n20196_not
g41880 not n14940 ; n14940_not
g41881 not n14823 ; n14823_not
g41882 not n10890 ; n10890_not
g41883 not n26901 ; n26901_not
g41884 not n26370 ; n26370_not
g41885 not n10755 ; n10755_not
g41886 not n16533 ; n16533_not
g41887 not n15606 ; n15606_not
g41888 not n10908 ; n10908_not
g41889 not n10557 ; n10557_not
g41890 not n26361 ; n26361_not
g41891 not n18126 ; n18126_not
g41892 not n24471 ; n24471_not
g41893 not n22644 ; n22644_not
g41894 not n24606 ; n24606_not
g41895 not n16713 ; n16713_not
g41896 not n23364 ; n23364_not
g41897 not n10917 ; n10917_not
g41898 not n10926 ; n10926_not
g41899 not n21429 ; n21429_not
g41900 not n26910 ; n26910_not
g41901 not n26352 ; n26352_not
g41902 not n15156 ; n15156_not
g41903 not n26433 ; n26433_not
g41904 not n22662 ; n22662_not
g41905 not n10872 ; n10872_not
g41906 not n18153 ; n18153_not
g41907 not n21636 ; n21636_not
g41908 not n24480 ; n24480_not
g41909 not n14832 ; n14832_not
g41910 not n26424 ; n26424_not
g41911 not n26325 ; n26325_not
g41912 not n23229 ; n23229_not
g41913 not n26415 ; n26415_not
g41914 not n22653 ; n22653_not
g41915 not n10566 ; n10566_not
g41916 not n23355 ; n23355_not
g41917 not n10881 ; n10881_not
g41918 not n18144 ; n18144_not
g41919 not n26343 ; n26343_not
g41920 not n14904 ; n14904_not
g41921 not n23256 ; n23256_not
g41922 not n10692 ; n10692_not
g41923 not n18306 ; n18306_not
g41924 not n26622 ; n26622_not
g41925 not n21825 ; n21825_not
g41926 not n23274 ; n23274_not
g41927 not n21654 ; n21654_not
g41928 not n26613 ; n26613_not
g41929 not n15534 ; n15534_not
g41930 not n24561 ; n24561_not
g41931 not n13554 ; n13554_not
g41932 not n10719 ; n10719_not
g41933 not n10638 ; n10638_not
g41934 not n22770 ; n22770_not
g41935 not n22761 ; n22761_not
g41936 not n16362 ; n16362_not
g41937 not n10737 ; n10737_not
g41938 not n26712 ; n26712_not
g41939 not n15507 ; n15507_not
g41940 not n14913 ; n14913_not
g41941 not n24552 ; n24552_not
g41942 not n10656 ; n10656_not
g41943 not n26703 ; n26703_not
g41944 not n10674 ; n10674_not
g41945 not n15516 ; n15516_not
g41946 not n14652 ; n14652_not
g41947 not n23265 ; n23265_not
g41948 not n21663 ; n21663_not
g41949 not n26721 ; n26721_not
g41950 not n15525 ; n15525_not
g41951 not n10683 ; n10683_not
g41952 not n26640 ; n26640_not
g41953 not n26631 ; n26631_not
g41954 not n22734 ; n22734_not
g41955 not n23292 ; n23292_not
g41956 not n26532 ; n26532_not
g41957 not n22806 ; n22806_not
g41958 not n10593 ; n10593_not
g41959 not n10782 ; n10782_not
g41960 not n18225 ; n18225_not
g41961 not n26523 ; n26523_not
g41962 not n21645 ; n21645_not
g41963 not n26514 ; n26514_not
g41964 not n22725 ; n22725_not
g41965 not n16542 ; n16542_not
g41966 not n18216 ; n18216_not
g41967 not n13383 ; n13383_not
g41968 not n23319 ; n23319_not
g41969 not n20178 ; n20178_not
g41970 not n20088 ; n20088_not
g41971 not n26811 ; n26811_not
g41972 not n18261 ; n18261_not
g41973 not n22752 ; n22752_not
g41974 not n24381 ; n24381_not
g41975 not n26604 ; n26604_not
g41976 not n10629 ; n10629_not
g41977 not n24570 ; n24570_not
g41978 not n20097 ; n20097_not
g41979 not n23283 ; n23283_not
g41980 not n22743 ; n22743_not
g41981 not n10539 ; n10539_not
g41982 not n14931 ; n14931_not
g41983 not n26730 ; n26730_not
g41984 not n10764 ; n10764_not
g41985 not n23247 ; n23247_not
g41986 not n18243 ; n18243_not
g41987 not n15552 ; n15552_not
g41988 not n18315 ; n18315_not
g41989 not n15543 ; n15543_not
g41990 not n10458 ; n10458_not
g41991 not n26550 ; n26550_not
g41992 not n26802 ; n26802_not
g41993 not n26235 ; n26235_not
g41994 not n22716 ; n22716_not
g41995 not n13347 ; n13347_not
g41996 not n22581 ; n22581_not
g41997 not n16524 ; n16524_not
g41998 not n21816 ; n21816_not
g41999 not n11259 ; n11259_not
g42000 not n15444 ; n15444_not
g42001 not n22563 ; n22563_not
g42002 not n11268 ; n11268_not
g42003 not n13338 ; n13338_not
g42004 not n26226 ; n26226_not
g42005 not n11286 ; n11286_not
g42006 not n13473 ; n13473_not
g42007 not n14733 ; n14733_not
g42008 not n13572 ; n13572_not
g42009 not n23463 ; n23463_not
g42010 not n22545 ; n22545_not
g42011 not n14292 ; n14292_not
g42012 not n24462 ; n24462_not
g42013 not n21609 ; n21609_not
g42014 not n23472 ; n23472_not
g42015 not n26244 ; n26244_not
g42016 not n14760 ; n14760_not
g42017 not n22860 ; n22860_not
g42018 not n24624 ; n24624_not
g42019 not n15228 ; n15228_not
g42020 not n23445 ; n23445_not
g42021 not n14751 ; n14751_not
g42022 not n11169 ; n11169_not
g42023 not n16731 ; n16731_not
g42024 not n11178 ; n11178_not
g42025 not n10368 ; n10368_not
g42026 not n23454 ; n23454_not
g42027 not n11187 ; n11187_not
g42028 not n10449 ; n10449_not
g42029 not n22590 ; n22590_not
g42030 not n11196 ; n11196_not
g42031 not n15264 ; n15264_not
g42032 not n14706 ; n14706_not
g42033 not n20367 ; n20367_not
g42034 not n10386 ; n10386_not
g42035 not n16515 ; n16515_not
g42036 not n11376 ; n11376_not
g42037 not n15714 ; n15714_not
g42038 not n23481 ; n23481_not
g42039 not n20376 ; n20376_not
g42040 not n22527 ; n22527_not
g42041 not n11385 ; n11385_not
g42042 not n10377 ; n10377_not
g42043 not n23490 ; n23490_not
g42044 not n20385 ; n20385_not
g42045 not n11394 ; n11394_not
g42046 not n23166 ; n23166_not
g42047 not n20394 ; n20394_not
g42048 not n27018 ; n27018_not
g42049 not n14724 ; n14724_not
g42050 not n23409 ; n23409_not
g42051 not n20349 ; n20349_not
g42052 not n16740 ; n16740_not
g42053 not n15705 ; n15705_not
g42054 not n14715 ; n14715_not
g42055 not n11358 ; n11358_not
g42056 not n11349 ; n11349_not
g42057 not n13545 ; n13545_not
g42058 not n10395 ; n10395_not
g42059 not n21852 ; n21852_not
g42060 not n26217 ; n26217_not
g42061 not n23175 ; n23175_not
g42062 not n22536 ; n22536_not
g42063 not n27306 ; n27306_not
g42064 not n10962 ; n10962_not
g42065 not n18090 ; n18090_not
g42066 not n26316 ; n26316_not
g42067 not n15174 ; n15174_not
g42068 not n10971 ; n10971_not
g42069 not n21681 ; n21681_not
g42070 not n23382 ; n23382_not
g42071 not n20268 ; n20268_not
g42072 not n18081 ; n18081_not
g42073 not n21690 ; n21690_not
g42074 not n26307 ; n26307_not
g42075 not n10980 ; n10980_not
g42076 not n18072 ; n18072_not
g42077 not n16407 ; n16407_not
g42078 not n20277 ; n20277_not
g42079 not n15462 ; n15462_not
g42080 not n14814 ; n14814_not
g42081 not n18117 ; n18117_not
g42082 not n10935 ; n10935_not
g42083 not n15471 ; n15471_not
g42084 not n23148 ; n23148_not
g42085 not n13365 ; n13365_not
g42086 not n14805 ; n14805_not
g42087 not n10944 ; n10944_not
g42088 not n26334 ; n26334_not
g42089 not n10953 ; n10953_not
g42090 not n24615 ; n24615_not
g42091 not n10548 ; n10548_not
g42092 not n15624 ; n15624_not
g42093 not n22833 ; n22833_not
g42094 not n18360 ; n18360_not
g42095 not n18045 ; n18045_not
g42096 not n12942 ; n12942_not
g42097 not n23418 ; n23418_not
g42098 not n10476 ; n10476_not
g42099 not n15651 ; n15651_not
g42100 not n11079 ; n11079_not
g42101 not n18036 ; n18036_not
g42102 not n14607 ; n14607_not
g42103 not n11097 ; n11097_not
g42104 not n10467 ; n10467_not
g42105 not n15660 ; n15660_not
g42106 not n18027 ; n18027_not
g42107 not n23436 ; n23436_not
g42108 not n23193 ; n23193_not
g42109 not n26271 ; n26271_not
g42110 not n21843 ; n21843_not
g42111 not n20286 ; n20286_not
g42112 not n18063 ; n18063_not
g42113 not n15642 ; n15642_not
g42114 not n26262 ; n26262_not
g42115 not n13356 ; n13356_not
g42116 not n13419 ; n13419_not
g42117 not n22851 ; n22851_not
g42118 not n20295 ; n20295_not
g42119 not n10728 ; n10728_not
g42120 not n18054 ; n18054_not
g42121 not n16722 ; n16722_not
g42122 not n10485 ; n10485_not
g42123 not n15453 ; n15453_not
g42124 not n26253 ; n26253_not
g42125 not n12573 ; n12573_not
g42126 not n13941 ; n13941_not
g42127 not n25308 ; n25308_not
g42128 not n12690 ; n12690_not
g42129 not n24804 ; n24804_not
g42130 not n12582 ; n12582_not
g42131 not n18630 ; n18630_not
g42132 not n25263 ; n25263_not
g42133 not n16425 ; n16425_not
g42134 not n25290 ; n25290_not
g42135 not n13932 ; n13932_not
g42136 not n19062 ; n19062_not
g42137 not n16605 ; n16605_not
g42138 not n12546 ; n12546_not
g42139 not n12609 ; n12609_not
g42140 not n27063 ; n27063_not
g42141 not n23076 ; n23076_not
g42142 not n25272 ; n25272_not
g42143 not n20916 ; n20916_not
g42144 not n16227 ; n16227_not
g42145 not n21366 ; n21366_not
g42146 not n13059 ; n13059_not
g42147 not n17226 ; n17226_not
g42148 not n16434 ; n16434_not
g42149 not n25326 ; n25326_not
g42150 not n24129 ; n24129_not
g42151 not n19071 ; n19071_not
g42152 not n16209 ; n16209_not
g42153 not n12555 ; n12555_not
g42154 not n24138 ; n24138_not
g42155 not n13950 ; n13950_not
g42156 not n24390 ; n24390_not
g42157 not n12564 ; n12564_not
g42158 not n17208 ; n17208_not
g42159 not n24714 ; n24714_not
g42160 not n23922 ; n23922_not
g42161 not n24147 ; n24147_not
g42162 not n16245 ; n16245_not
g42163 not n12654 ; n12654_not
g42164 not n24174 ; n24174_not
g42165 not n27180 ; n27180_not
g42166 not n16236 ; n16236_not
g42167 not n16902 ; n16902_not
g42168 not n24183 ; n24183_not
g42169 not n21195 ; n21195_not
g42170 not n27090 ; n27090_not
g42171 not n17154 ; n17154_not
g42172 not n12672 ; n12672_not
g42173 not n24831 ; n24831_not
g42174 not n16074 ; n16074_not
g42175 not n25236 ; n25236_not
g42176 not n17145 ; n17145_not
g42177 not n13860 ; n13860_not
g42178 not n24840 ; n24840_not
g42179 not n25227 ; n25227_not
g42180 not n19035 ; n19035_not
g42181 not n17190 ; n17190_not
g42182 not n24156 ; n24156_not
g42183 not n12627 ; n12627_not
g42184 not n13923 ; n13923_not
g42185 not n18720 ; n18720_not
g42186 not n13671 ; n13671_not
g42187 not n24165 ; n24165_not
g42188 not n19044 ; n19044_not
g42189 not n12636 ; n12636_not
g42190 not n27153 ; n27153_not
g42191 not n13914 ; n13914_not
g42192 not n25254 ; n25254_not
g42193 not n17172 ; n17172_not
g42194 not n24822 ; n24822_not
g42195 not n13905 ; n13905_not
g42196 not n17163 ; n17163_not
g42197 not n19107 ; n19107_not
g42198 not n22158 ; n22158_not
g42199 not n12438 ; n12438_not
g42200 not n12447 ; n12447_not
g42201 not n14076 ; n14076_not
g42202 not n12456 ; n12456_not
g42203 not n22167 ; n22167_not
g42204 not n13086 ; n13086_not
g42205 not n25380 ; n25380_not
g42206 not n17280 ; n17280_not
g42207 not n25371 ; n25371_not
g42208 not n15237 ; n15237_not
g42209 not n18621 ; n18621_not
g42210 not n27081 ; n27081_not
g42211 not n24075 ; n24075_not
g42212 not n17271 ; n17271_not
g42213 not n14067 ; n14067_not
g42214 not n12474 ; n12474_not
g42215 not n21438 ; n21438_not
g42216 not n25362 ; n25362_not
g42217 not n16443 ; n16443_not
g42218 not n17316 ; n17316_not
g42219 not n12375 ; n12375_not
g42220 not n27072 ; n27072_not
g42221 not n24732 ; n24732_not
g42222 not n27207 ; n27207_not
g42223 not n25416 ; n25416_not
g42224 not n24057 ; n24057_not
g42225 not n25317 ; n25317_not
g42226 not n14094 ; n14094_not
g42227 not n12393 ; n12393_not
g42228 not n24066 ; n24066_not
g42229 not n13482 ; n13482_not
g42230 not n14085 ; n14085_not
g42231 not n12339 ; n12339_not
g42232 not n24750 ; n24750_not
g42233 not n16137 ; n16137_not
g42234 not n21771 ; n21771_not
g42235 not n12429 ; n12429_not
g42236 not n21159 ; n21159_not
g42237 not n21942 ; n21942_not
g42238 not n24084 ; n24084_not
g42239 not n13068 ; n13068_not
g42240 not n16182 ; n16182_not
g42241 not n17244 ; n17244_not
g42242 not n12519 ; n12519_not
g42243 not n22149 ; n22149_not
g42244 not n19080 ; n19080_not
g42245 not n21168 ; n21168_not
g42246 not n12528 ; n12528_not
g42247 not n13662 ; n13662_not
g42248 not n16191 ; n16191_not
g42249 not n17235 ; n17235_not
g42250 not n15318 ; n15318_not
g42251 not n24093 ; n24093_not
g42252 not n25335 ; n25335_not
g42253 not n21177 ; n21177_not
g42254 not n25218 ; n25218_not
g42255 not n16146 ; n16146_not
g42256 not n16155 ; n16155_not
g42257 not n14058 ; n14058_not
g42258 not n25353 ; n25353_not
g42259 not n24408 ; n24408_not
g42260 not n12483 ; n12483_not
g42261 not n14049 ; n14049_not
g42262 not n16164 ; n16164_not
g42263 not n12492 ; n12492_not
g42264 not n13653 ; n13653_not
g42265 not n18612 ; n18612_not
g42266 not n17253 ; n17253_not
g42267 not n25344 ; n25344_not
g42268 not n24363 ; n24363_not
g42269 not n12843 ; n12843_not
g42270 not n24309 ; n24309_not
g42271 not n12618 ; n12618_not
g42272 not n22068 ; n22068_not
g42273 not n17019 ; n17019_not
g42274 not n12852 ; n12852_not
g42275 not n24354 ; n24354_not
g42276 not n18900 ; n18900_not
g42277 not n25092 ; n25092_not
g42278 not n16353 ; n16353_not
g42279 not n13761 ; n13761_not
g42280 not n24255 ; n24255_not
g42281 not n24318 ; n24318_not
g42282 not n18810 ; n18810_not
g42283 not n13752 ; n13752_not
g42284 not n24912 ; n24912_not
g42285 not n12870 ; n12870_not
g42286 not n25074 ; n25074_not
g42287 not n25119 ; n25119_not
g42288 not n21285 ; n21285_not
g42289 not n21276 ; n21276_not
g42290 not n17046 ; n17046_not
g42291 not n23058 ; n23058_not
g42292 not n12816 ; n12816_not
g42293 not n13680 ; n13680_not
g42294 not n24282 ; n24282_not
g42295 not n27135 ; n27135_not
g42296 not n24291 ; n24291_not
g42297 not n12825 ; n12825_not
g42298 not n17037 ; n17037_not
g42299 not n12834 ; n12834_not
g42300 not n24507 ; n24507_not
g42301 not n13770 ; n13770_not
g42302 not n21294 ; n21294_not
g42303 not n24903 ; n24903_not
g42304 not n21375 ; n21375_not
g42305 not n16344 ; n16344_not
g42306 not n27126 ; n27126_not
g42307 not n16380 ; n16380_not
g42308 not n12591 ; n12591_not
g42309 not n13725 ; n13725_not
g42310 not n12933 ; n12933_not
g42311 not n25029 ; n25029_not
g42312 not n21339 ; n21339_not
g42313 not n24336 ; n24336_not
g42314 not n13716 ; n13716_not
g42315 not n21357 ; n21357_not
g42316 not n18702 ; n18702_not
g42317 not n24345 ; n24345_not
g42318 not n12951 ; n12951_not
g42319 not n15282 ; n15282_not
g42320 not n21348 ; n21348_not
g42321 not n13509 ; n13509_not
g42322 not n12960 ; n12960_not
g42323 not n25065 ; n25065_not
g42324 not n18801 ; n18801_not
g42325 not n25056 ; n25056_not
g42326 not n24327 ; n24327_not
g42327 not n16470 ; n16470_not
g42328 not n25047 ; n25047_not
g42329 not n18531 ; n18531_not
g42330 not n25038 ; n25038_not
g42331 not n13743 ; n13743_not
g42332 not n16371 ; n16371_not
g42333 not n13734 ; n13734_not
g42334 not n24930 ; n24930_not
g42335 not n12915 ; n12915_not
g42336 not n12906 ; n12906_not
g42337 not n21753 ; n21753_not
g42338 not n12924 ; n12924_not
g42339 not n21249 ; n21249_not
g42340 not n27162 ; n27162_not
g42341 not n17118 ; n17118_not
g42342 not n22095 ; n22095_not
g42343 not n12726 ; n12726_not
g42344 not n17109 ; n17109_not
g42345 not n16290 ; n16290_not
g42346 not n25209 ; n25209_not
g42347 not n13824 ; n13824_not
g42348 not n19026 ; n19026_not
g42349 not n27045 ; n27045_not
g42350 not n12735 ; n12735_not
g42351 not n12744 ; n12744_not
g42352 not n15255 ; n15255_not
g42353 not n15309 ; n15309_not
g42354 not n25182 ; n25182_not
g42355 not n22086 ; n22086_not
g42356 not n12753 ; n12753_not
g42357 not n19017 ; n19017_not
g42358 not n13815 ; n13815_not
g42359 not n12681 ; n12681_not
g42360 not n12645 ; n12645_not
g42361 not n17127 ; n17127_not
g42362 not n17136 ; n17136_not
g42363 not n13851 ; n13851_not
g42364 not n24219 ; n24219_not
g42365 not n16272 ; n16272_not
g42366 not n13842 ; n13842_not
g42367 not n21393 ; n21393_not
g42368 not n24372 ; n24372_not
g42369 not n12708 ; n12708_not
g42370 not n24228 ; n24228_not
g42371 not n27171 ; n27171_not
g42372 not n21762 ; n21762_not
g42373 not n17028 ; n17028_not
g42374 not n24264 ; n24264_not
g42375 not n13491 ; n13491_not
g42376 not n21384 ; n21384_not
g42377 not n25137 ; n25137_not
g42378 not n16317 ; n16317_not
g42379 not n16920 ; n16920_not
g42380 not n27108 ; n27108_not
g42381 not n25128 ; n25128_not
g42382 not n17064 ; n17064_not
g42383 not n16416 ; n16416_not
g42384 not n17055 ; n17055_not
g42385 not n16326 ; n16326_not
g42386 not n22077 ; n22077_not
g42387 not n12807 ; n12807_not
g42388 not n15273 ; n15273_not
g42389 not n21744 ; n21744_not
g42390 not n24246 ; n24246_not
g42391 not n25164 ; n25164_not
g42392 not n21258 ; n21258_not
g42393 not n17091 ; n17091_not
g42394 not n16911 ; n16911_not
g42395 not n17082 ; n17082_not
g42396 not n12771 ; n12771_not
g42397 not n16308 ; n16308_not
g42398 not n21267 ; n21267_not
g42399 not n27144 ; n27144_not
g42400 not n25146 ; n25146_not
g42401 not n23067 ; n23067_not
g42402 not n21735 ; n21735_not
g42403 not n17505 ; n17505_not
g42404 not n16623 ; n16623_not
g42405 not n27261 ; n27261_not
g42406 not n23850 ; n23850_not
g42407 not n25425 ; n25425_not
g42408 not n20925 ; n20925_not
g42409 not n14364 ; n14364_not
g42410 not n27252 ; n27252_not
g42411 not n15165 ; n15165_not
g42412 not n21780 ; n21780_not
g42413 not n21492 ; n21492_not
g42414 not n25560 ; n25560_not
g42415 not n24705 ; n24705_not
g42416 not n21933 ; n21933_not
g42417 not n20907 ; n20907_not
g42418 not n17523 ; n17523_not
g42419 not n11961 ; n11961_not
g42420 not n19242 ; n19242_not
g42421 not n27270 ; n27270_not
g42422 not n25623 ; n25623_not
g42423 not n23832 ; n23832_not
g42424 not n14382 ; n14382_not
g42425 not n15147 ; n15147_not
g42426 not n19224 ; n19224_not
g42427 not n13185 ; n13185_not
g42428 not n23841 ; n23841_not
g42429 not n14373 ; n14373_not
g42430 not n19170 ; n19170_not
g42431 not n17460 ; n17460_not
g42432 not n23904 ; n23904_not
g42433 not n11853 ; n11853_not
g42434 not n24426 ; n24426_not
g42435 not n14328 ; n14328_not
g42436 not n14319 ; n14319_not
g42437 not n24417 ; n24417_not
g42438 not n13635 ; n13635_not
g42439 not n12078 ; n12078_not
g42440 not n23913 ; n23913_not
g42441 not n19152 ; n19152_not
g42442 not n25524 ; n25524_not
g42443 not n17442 ; n17442_not
g42444 not n20934 ; n20934_not
g42445 not n15345 ; n15345_not
g42446 not n24525 ; n24525_not
g42447 not n25551 ; n25551_not
g42448 not n14355 ; n14355_not
g42449 not n20952 ; n20952_not
g42450 not n27243 ; n27243_not
g42451 not n25542 ; n25542_not
g42452 not n13626 ; n13626_not
g42453 not n14346 ; n14346_not
g42454 not n20970 ; n20970_not
g42455 not n27054 ; n27054_not
g42456 not n14337 ; n14337_not
g42457 not n25533 ; n25533_not
g42458 not n16830 ; n16830_not
g42459 not n11907 ; n11907_not
g42460 not n10098 ; n10098_not
g42461 not n22275 ; n22275_not
g42462 not n20808 ; n20808_not
g42463 not n11916 ; n11916_not
g42464 not n19332 ; n19332_not
g42465 not n25740 ; n25740_not
g42466 not n19323 ; n19323_not
g42467 not n19314 ; n19314_not
g42468 not n18405 ; n18405_not
g42469 not n25731 ; n25731_not
g42470 not n14427 ; n14427_not
g42471 not n16812 ; n16812_not
g42472 not n20817 ; n20817_not
g42473 not n11925 ; n11925_not
g42474 not n11934 ; n11934_not
g42475 not n25722 ; n25722_not
g42476 not n20628 ; n20628_not
g42477 not n25803 ; n25803_not
g42478 not n23805 ; n23805_not
g42479 not n19350 ; n19350_not
g42480 not n20763 ; n20763_not
g42481 not n15093 ; n15093_not
g42482 not n21519 ; n21519_not
g42483 not n16632 ; n16632_not
g42484 not n14436 ; n14436_not
g42485 not n22941 ; n22941_not
g42486 not n20781 ; n20781_not
g42487 not n22284 ; n22284_not
g42488 not n20790 ; n20790_not
g42489 not n25704 ; n25704_not
g42490 not n20853 ; n20853_not
g42491 not n15129 ; n15129_not
g42492 not n11880 ; n11880_not
g42493 not n23814 ; n23814_not
g42494 not n15066 ; n15066_not
g42495 not n20862 ; n20862_not
g42496 not n11952 ; n11952_not
g42497 not n22248 ; n22248_not
g42498 not n20871 ; n20871_not
g42499 not n20880 ; n20880_not
g42500 not n17532 ; n17532_not
g42501 not n25650 ; n25650_not
g42502 not n19260 ; n19260_not
g42503 not n25632 ; n25632_not
g42504 not n14418 ; n14418_not
g42505 not n25713 ; n25713_not
g42506 not n10089 ; n10089_not
g42507 not n20826 ; n20826_not
g42508 not n15363 ; n15363_not
g42509 not n20835 ; n20835_not
g42510 not n14409 ; n14409_not
g42511 not n13077 ; n13077_not
g42512 not n11943 ; n11943_not
g42513 not n20844 ; n20844_not
g42514 not n14391 ; n14391_not
g42515 not n17550 ; n17550_not
g42516 not n19305 ; n19305_not
g42517 not n12348 ; n12348_not
g42518 not n13158 ; n13158_not
g42519 not n13149 ; n13149_not
g42520 not n22176 ; n22176_not
g42521 not n21087 ; n21087_not
g42522 not n12177 ; n12177_not
g42523 not n14229 ; n14229_not
g42524 not n14175 ; n14175_not
g42525 not n19116 ; n19116_not
g42526 not n19134 ; n19134_not
g42527 not n16452 ; n16452_not
g42528 not n14256 ; n14256_not
g42529 not n18351 ; n18351_not
g42530 not n12186 ; n12186_not
g42531 not n25434 ; n25434_not
g42532 not n14166 ; n14166_not
g42533 not n13518 ; n13518_not
g42534 not n25506 ; n25506_not
g42535 not n17343 ; n17343_not
g42536 not n14247 ; n14247_not
g42537 not n27225 ; n27225_not
g42538 not n12195 ; n12195_not
g42539 not n14238 ; n14238_not
g42540 not n17361 ; n17361_not
g42541 not n12276 ; n12276_not
g42542 not n13806 ; n13806_not
g42543 not n25443 ; n25443_not
g42544 not n17370 ; n17370_not
g42545 not n23085 ; n23085_not
g42546 not n12285 ; n12285_not
g42547 not n14184 ; n14184_not
g42548 not n12294 ; n12294_not
g42549 not n25470 ; n25470_not
g42550 not n25461 ; n25461_not
g42551 not n19125 ; n19125_not
g42552 not n12717 ; n12717_not
g42553 not n25452 ; n25452_not
g42554 not n23094 ; n23094_not
g42555 not n12249 ; n12249_not
g42556 not n21924 ; n21924_not
g42557 not n15192 ; n15192_not
g42558 not n21456 ; n21456_not
g42559 not n21960 ; n21960_not
g42560 not n21069 ; n21069_not
g42561 not n12267 ; n12267_not
g42562 not n16614 ; n16614_not
g42563 not n16083 ; n16083_not
g42564 not n21078 ; n21078_not
g42565 not n24723 ; n24723_not
g42566 not n12159 ; n12159_not
g42567 not n27216 ; n27216_not
g42568 not n21951 ; n21951_not
g42569 not n14274 ; n14274_not
g42570 not n13095 ; n13095_not
g42571 not n16119 ; n16119_not
g42572 not n14283 ; n14283_not
g42573 not n12366 ; n12366_not
g42574 not n23940 ; n23940_not
g42575 not n13644 ; n13644_not
g42576 not n15183 ; n15183_not
g42577 not n14139 ; n14139_not
g42578 not n13833 ; n13833_not
g42579 not n23931 ; n23931_not
g42580 not n17433 ; n17433_not
g42581 not n12096 ; n12096_not
g42582 not n21483 ; n21483_not
g42583 not n16038 ; n16038_not
g42584 not n13167 ; n13167_not
g42585 not n24048 ; n24048_not
g42586 not n12168 ; n12168_not
g42587 not n14148 ; n14148_not
g42588 not n21096 ; n21096_not
g42589 not n21474 ; n21474_not
g42590 not n17415 ; n17415_not
g42591 not n12357 ; n12357_not
g42592 not n23823 ; n23823_not
g42593 not n14265 ; n14265_not
g42594 not n16056 ; n16056_not
g42595 not n24039 ; n24039_not
g42596 not n19063 ; n19063_not
g42597 not n27217 ; n27217_not
g42598 not n18730 ; n18730_not
g42599 not n24535 ; n24535_not
g42600 not n21790 ; n21790_not
g42601 not n19306 ; n19306_not
g42602 not n23239 ; n23239_not
g42603 not n27073 ; n27073_not
g42604 not n20089 ; n20089_not
g42605 not n18604 ; n18604_not
g42606 not n21754 ; n21754_not
g42607 not n19423 ; n19423_not
g42608 not n19333 ; n19333_not
g42609 not n26812 ; n26812_not
g42610 not n27136 ; n27136_not
g42611 not n27037 ; n27037_not
g42612 not n19108 ; n19108_not
g42613 not n22771 ; n22771_not
g42614 not n19630 ; n19630_not
g42615 not n19360 ; n19360_not
g42616 not n19324 ; n19324_not
g42617 not n23086 ; n23086_not
g42618 not n19351 ; n19351_not
g42619 not n18541 ; n18541_not
g42620 not n18505 ; n18505_not
g42621 not n27190 ; n27190_not
g42622 not n21772 ; n21772_not
g42623 not n24364 ; n24364_not
g42624 not n18811 ; n18811_not
g42625 not n19405 ; n19405_not
g42626 not n23257 ; n23257_not
g42627 not n26722 ; n26722_not
g42628 not n23158 ; n23158_not
g42629 not n27028 ; n27028_not
g42630 not n26713 ; n26713_not
g42631 not n26731 ; n26731_not
g42632 not n18802 ; n18802_not
g42633 not n23248 ; n23248_not
g42634 not n21628 ; n21628_not
g42635 not n21745 ; n21745_not
g42636 not n18910 ; n18910_not
g42637 not n21727 ; n21727_not
g42638 not n22807 ; n22807_not
g42639 not n19018 ; n19018_not
g42640 not n18703 ; n18703_not
g42641 not n27208 ; n27208_not
g42642 not n18712 ; n18712_not
g42643 not n19315 ; n19315_not
g42644 not n22906 ; n22906_not
g42645 not n19117 ; n19117_not
g42646 not n21673 ; n21673_not
g42647 not n18820 ; n18820_not
g42648 not n21808 ; n21808_not
g42649 not n26803 ; n26803_not
g42650 not n27127 ; n27127_not
g42651 not n23167 ; n23167_not
g42652 not n27055 ; n27055_not
g42653 not n19414 ; n19414_not
g42654 not n19441 ; n19441_not
g42655 not n19036 ; n19036_not
g42656 not n26911 ; n26911_not
g42657 not n19540 ; n19540_not
g42658 not n19531 ; n19531_not
g42659 not n23194 ; n23194_not
g42660 not n22915 ; n22915_not
g42661 not n27091 ; n27091_not
g42662 not n19522 ; n19522_not
g42663 not n27244 ; n27244_not
g42664 not n23176 ; n23176_not
g42665 not n21718 ; n21718_not
g42666 not n19513 ; n19513_not
g42667 not n27226 ; n27226_not
g42668 not n19207 ; n19207_not
g42669 not n19504 ; n19504_not
g42670 not n22870 ; n22870_not
g42671 not n19027 ; n19027_not
g42672 not n19072 ; n19072_not
g42673 not n27253 ; n27253_not
g42674 not n19045 ; n19045_not
g42675 not n22852 ; n22852_not
g42676 not n27181 ; n27181_not
g42677 not n21817 ; n21817_not
g42678 not n26902 ; n26902_not
g42679 not n26920 ; n26920_not
g42680 not n21763 ; n21763_not
g42681 not n19342 ; n19342_not
g42682 not n24490 ; n24490_not
g42683 not n19612 ; n19612_not
g42684 not n19621 ; n19621_not
g42685 not n19153 ; n19153_not
g42686 not n19603 ; n19603_not
g42687 not n19144 ; n19144_not
g42688 not n19801 ; n19801_not
g42689 not n21691 ; n21691_not
g42690 not n27235 ; n27235_not
g42691 not n23095 ; n23095_not
g42692 not n27172 ; n27172_not
g42693 not n19135 ; n19135_not
g42694 not n19171 ; n19171_not
g42695 not n22834 ; n22834_not
g42696 not n21781 ; n21781_not
g42697 not n26821 ; n26821_not
g42698 not n19090 ; n19090_not
g42699 not n19081 ; n19081_not
g42700 not n23185 ; n23185_not
g42701 not n24544 ; n24544_not
g42702 not n27307 ; n27307_not
g42703 not n19243 ; n19243_not
g42704 not n19252 ; n19252_not
g42705 not n27064 ; n27064_not
g42706 not n22951 ; n22951_not
g42707 not n24508 ; n24508_not
g42708 not n19720 ; n19720_not
g42709 not n19261 ; n19261_not
g42710 not n22564 ; n22564_not
g42711 not n27109 ; n27109_not
g42712 not n22465 ; n22465_not
g42713 not n19900 ; n19900_not
g42714 not n19126 ; n19126_not
g42715 not n27271 ; n27271_not
g42716 not n27046 ; n27046_not
g42717 not n23059 ; n23059_not
g42718 not n27019 ; n27019_not
g42719 not n24526 ; n24526_not
g42720 not n22924 ; n22924_not
g42721 not n27262 ; n27262_not
g42722 not n19702 ; n19702_not
g42723 not n22933 ; n22933_not
g42724 not n24517 ; n24517_not
g42725 not n22825 ; n22825_not
g42726 not n27163 ; n27163_not
g42727 not n27154 ; n27154_not
g42728 not n19450 ; n19450_not
g42729 not n19225 ; n19225_not
g42730 not n19711 ; n19711_not
g42731 not n21736 ; n21736_not
g42732 not n23077 ; n23077_not
g42733 not n22942 ; n22942_not
g42734 not n27145 ; n27145_not
g42735 not n22816 ; n22816_not
g42736 not n26830 ; n26830_not
g42737 not n25354 ; n25354_not
g42738 not n25534 ; n25534_not
g42739 not n20890 ; n20890_not
g42740 not n20971 ; n20971_not
g42741 not n20953 ; n20953_not
g42742 not n21934 ; n21934_not
g42743 not n20944 ; n20944_not
g42744 not n25552 ; n25552_not
g42745 not n25543 ; n25543_not
g42746 not n20935 ; n20935_not
g42747 not n25561 ; n25561_not
g42748 not n25462 ; n25462_not
g42749 not n25570 ; n25570_not
g42750 not n20926 ; n20926_not
g42751 not n23860 ; n23860_not
g42752 not n20917 ; n20917_not
g42753 not n23851 ; n23851_not
g42754 not n23662 ; n23662_not
g42755 not n25606 ; n25606_not
g42756 not n23842 ; n23842_not
g42757 not n23833 ; n23833_not
g42758 not n25615 ; n25615_not
g42759 not n24706 ; n24706_not
g42760 not n25624 ; n25624_not
g42761 not n25435 ; n25435_not
g42762 not n21079 ; n21079_not
g42763 not n22177 ; n22177_not
g42764 not n21457 ; n21457_not
g42765 not n22168 ; n22168_not
g42766 not n25444 ; n25444_not
g42767 not n25453 ; n25453_not
g42768 not n25408 ; n25408_not
g42769 not n25471 ; n25471_not
g42770 not n22186 ; n22186_not
g42771 not n21943 ; n21943_not
g42772 not n21466 ; n21466_not
g42773 not n22195 ; n22195_not
g42774 not n21952 ; n21952_not
g42775 not n21295 ; n21295_not
g42776 not n24715 ; n24715_not
g42777 not n21268 ; n21268_not
g42778 not n25507 ; n25507_not
g42779 not n21475 ; n21475_not
g42780 not n23824 ; n23824_not
g42781 not n23950 ; n23950_not
g42782 not n23941 ; n23941_not
g42783 not n23932 ; n23932_not
g42784 not n25516 ; n25516_not
g42785 not n23923 ; n23923_not
g42786 not n25525 ; n25525_not
g42787 not n21493 ; n21493_not
g42788 not n23905 ; n23905_not
g42789 not n20809 ; n20809_not
g42790 not n22276 ; n22276_not
g42791 not n25750 ; n25750_not
g42792 not n23806 ; n23806_not
g42793 not n20782 ; n20782_not
g42794 not n22285 ; n22285_not
g42795 not n21916 ; n21916_not
g42796 not n20764 ; n20764_not
g42797 not n22294 ; n22294_not
g42798 not n25804 ; n25804_not
g42799 not n20755 ; n20755_not
g42800 not n25813 ; n25813_not
g42801 not n23770 ; n23770_not
g42802 not n23761 ; n23761_not
g42803 not n20746 ; n20746_not
g42804 not n25822 ; n25822_not
g42805 not n23752 ; n23752_not
g42806 not n25831 ; n25831_not
g42807 not n25723 ; n25723_not
g42808 not n20737 ; n20737_not
g42809 not n20728 ; n20728_not
g42810 not n25903 ; n25903_not
g42811 not n24661 ; n24661_not
g42812 not n25921 ; n25921_not
g42813 not n25930 ; n25930_not
g42814 not n23743 ; n23743_not
g42815 not n20719 ; n20719_not
g42816 not n25912 ; n25912_not
g42817 not n20908 ; n20908_not
g42818 not n25633 ; n25633_not
g42819 not n21925 ; n21925_not
g42820 not n25651 ; n25651_not
g42821 not n20881 ; n20881_not
g42822 not n25660 ; n25660_not
g42823 not n20872 ; n20872_not
g42824 not n22249 ; n22249_not
g42825 not n23815 ; n23815_not
g42826 not n20854 ; n20854_not
g42827 not n20845 ; n20845_not
g42828 not n24670 ; n24670_not
g42829 not n20827 ; n20827_not
g42830 not n20836 ; n20836_not
g42831 not n25705 ; n25705_not
g42832 not n20566 ; n20566_not
g42833 not n22267 ; n22267_not
g42834 not n20818 ; n20818_not
g42835 not n25732 ; n25732_not
g42836 not n25741 ; n25741_not
g42837 not n24283 ; n24283_not
g42838 not n24274 ; n24274_not
g42839 not n21286 ; n21286_not
g42840 not n22078 ; n22078_not
g42841 not n24265 ; n24265_not
g42842 not n21277 ; n21277_not
g42843 not n25138 ; n25138_not
g42844 not n25147 ; n25147_not
g42845 not n21385 ; n21385_not
g42846 not n21259 ; n21259_not
g42847 not n25165 ; n25165_not
g42848 not n25174 ; n25174_not
g42849 not n24247 ; n24247_not
g42850 not n24157 ; n24157_not
g42851 not n22087 ; n22087_not
g42852 not n25183 ; n25183_not
g42853 not n24238 ; n24238_not
g42854 not n24652 ; n24652_not
g42855 not n24850 ; n24850_not
g42856 not n24175 ; n24175_not
g42857 not n21844 ; n21844_not
g42858 not n24841 ; n24841_not
g42859 not n22096 ; n22096_not
g42860 not n24229 ; n24229_not
g42861 not n21394 ; n21394_not
g42862 not n24256 ; n24256_not
g42863 not n24346 ; n24346_not
g42864 not n21349 ; n21349_not
g42865 not n21358 ; n21358_not
g42866 not n24337 ; n24337_not
g42867 not n24904 ; n24904_not
g42868 not n24931 ; n24931_not
g42869 not n24328 ; n24328_not
g42870 not n24922 ; n24922_not
g42871 not n25039 ; n25039_not
g42872 not n25048 ; n25048_not
g42873 not n25057 ; n25057_not
g42874 not n24913 ; n24913_not
g42875 not n25066 ; n25066_not
g42876 not n21367 ; n21367_not
g42877 not n25075 ; n25075_not
g42878 not n24355 ; n24355_not
g42879 not n25084 ; n25084_not
g42880 not n25093 ; n25093_not
g42881 not n22069 ; n22069_not
g42882 not n24292 ; n24292_not
g42883 not n21826 ; n21826_not
g42884 not n24085 ; n24085_not
g42885 not n25336 ; n25336_not
g42886 not n24751 ; n24751_not
g42887 not n25345 ; n25345_not
g42888 not n22159 ; n22159_not
g42889 not n21439 ; n21439_not
g42890 not n25363 ; n25363_not
g42891 not n25381 ; n25381_not
g42892 not n24076 ; n24076_not
g42893 not n21097 ; n21097_not
g42894 not n24742 ; n24742_not
g42895 not n24733 ; n24733_not
g42896 not n25417 ; n25417_not
g42897 not n24049 ; n24049_not
g42898 not n24409 ; n24409_not
g42899 not n21448 ; n21448_not
g42900 not n24724 ; n24724_not
g42901 not n21088 ; n21088_not
g42902 not n21970 ; n21970_not
g42903 not n25219 ; n25219_not
g42904 not n25228 ; n25228_not
g42905 not n24832 ; n24832_not
g42906 not n25237 ; n25237_not
g42907 not n24184 ; n24184_not
g42908 not n25246 ; n25246_not
g42909 not n24823 ; n24823_not
g42910 not n24382 ; n24382_not
g42911 not n25255 ; n25255_not
g42912 not n24166 ; n24166_not
g42913 not n24805 ; n24805_not
g42914 not n25273 ; n25273_not
g42915 not n25264 ; n25264_not
g42916 not n21196 ; n21196_not
g42917 not n25282 ; n25282_not
g42918 not n24148 ; n24148_not
g42919 not n24139 ; n24139_not
g42920 not n25318 ; n25318_not
g42921 not n24391 ; n24391_not
g42922 not n25327 ; n25327_not
g42923 not n21178 ; n21178_not
g42924 not n21169 ; n21169_not
g42925 not n24067 ; n24067_not
g42926 not n23392 ; n23392_not
g42927 not n26272 ; n26272_not
g42928 not n23383 ; n23383_not
g42929 not n26281 ; n26281_not
g42930 not n26209 ; n26209_not
g42931 not n26290 ; n26290_not
g42932 not n26308 ; n26308_not
g42933 not n20269 ; n20269_not
g42934 not n23374 ; n23374_not
g42935 not n26317 ; n26317_not
g42936 not n22636 ; n22636_not
g42937 not n23347 ; n23347_not
g42938 not n26326 ; n26326_not
g42939 not n26335 ; n26335_not
g42940 not n26344 ; n26344_not
g42941 not n23149 ; n23149_not
g42942 not n24607 ; n24607_not
g42943 not n26353 ; n26353_not
g42944 not n23365 ; n23365_not
g42945 not n26362 ; n26362_not
g42946 not n24472 ; n24472_not
g42947 not n26371 ; n26371_not
g42948 not n26380 ; n26380_not
g42949 not n23356 ; n23356_not
g42950 not n22645 ; n22645_not
g42951 not n23473 ; n23473_not
g42952 not n22546 ; n22546_not
g42953 not n26227 ; n26227_not
g42954 not n22555 ; n22555_not
g42955 not n21619 ; n21619_not
g42956 not n22573 ; n22573_not
g42957 not n27316 ; n27316_not
g42958 not n26236 ; n26236_not
g42959 not n22582 ; n22582_not
g42960 not n23455 ; n23455_not
g42961 not n22591 ; n22591_not
g42962 not n22366 ; n22366_not
g42963 not n22609 ; n22609_not
g42964 not n23437 ; n23437_not
g42965 not n26245 ; n26245_not
g42966 not n23428 ; n23428_not
g42967 not n23419 ; n23419_not
g42968 not n22618 ; n22618_not
g42969 not n24463 ; n24463_not
g42970 not n20296 ; n20296_not
g42971 not n26254 ; n26254_not
g42972 not n20287 ; n20287_not
g42973 not n20197 ; n20197_not
g42974 not n23293 ; n23293_not
g42975 not n22735 ; n22735_not
g42976 not n26542 ; n26542_not
g42977 not n26551 ; n26551_not
g42978 not n24580 ; n24580_not
g42979 not n21646 ; n21646_not
g42980 not n23284 ; n23284_not
g42981 not n24481 ; n24481_not
g42982 not n26560 ; n26560_not
g42983 not n24571 ; n24571_not
g42984 not n26515 ; n26515_not
g42985 not n26605 ; n26605_not
g42986 not n22753 ; n22753_not
g42987 not n24562 ; n24562_not
g42988 not n23275 ; n23275_not
g42989 not n26623 ; n26623_not
g42990 not n26614 ; n26614_not
g42991 not n22780 ; n22780_not
g42992 not n26641 ; n26641_not
g42993 not n21664 ; n21664_not
g42994 not n26704 ; n26704_not
g42995 not n22654 ; n22654_not
g42996 not n26416 ; n26416_not
g42997 not n26425 ; n26425_not
g42998 not n26434 ; n26434_not
g42999 not n22663 ; n22663_not
g43000 not n21637 ; n21637_not
g43001 not n26443 ; n26443_not
g43002 not n26407 ; n26407_not
g43003 not n21835 ; n21835_not
g43004 not n26452 ; n26452_not
g43005 not n22672 ; n22672_not
g43006 not n26470 ; n26470_not
g43007 not n22681 ; n22681_not
g43008 not n22690 ; n22690_not
g43009 not n23338 ; n23338_not
g43010 not n26506 ; n26506_not
g43011 not n22717 ; n22717_not
g43012 not n20179 ; n20179_not
g43013 not n22726 ; n22726_not
g43014 not n26524 ; n26524_not
g43015 not n20494 ; n20494_not
g43016 not n21880 ; n21880_not
g43017 not n22384 ; n22384_not
g43018 not n22393 ; n22393_not
g43019 not n21709 ; n21709_not
g43020 not n20593 ; n20593_not
g43021 not n23653 ; n23653_not
g43022 not n23644 ; n23644_not
g43023 not n26083 ; n26083_not
g43024 not n20575 ; n20575_not
g43025 not n24643 ; n24643_not
g43026 not n21484 ; n21484_not
g43027 not n26074 ; n26074_not
g43028 not n21547 ; n21547_not
g43029 not n23635 ; n23635_not
g43030 not n26092 ; n26092_not
g43031 not n20548 ; n20548_not
g43032 not n21871 ; n21871_not
g43033 not n23617 ; n23617_not
g43034 not n26119 ; n26119_not
g43035 not n24436 ; n24436_not
g43036 not n23734 ; n23734_not
g43037 not n20665 ; n20665_not
g43038 not n23725 ; n23725_not
g43039 not n20683 ; n20683_not
g43040 not n20692 ; n20692_not
g43041 not n22339 ; n22339_not
g43042 not n21529 ; n21529_not
g43043 not n20674 ; n20674_not
g43044 not n23716 ; n23716_not
g43045 not n23707 ; n23707_not
g43046 not n22348 ; n22348_not
g43047 not n26029 ; n26029_not
g43048 not n20647 ; n20647_not
g43049 not n26038 ; n26038_not
g43050 not n20638 ; n20638_not
g43051 not n22357 ; n22357_not
g43052 not n20629 ; n20629_not
g43053 not n23680 ; n23680_not
g43054 not n20449 ; n20449_not
g43055 not n26056 ; n26056_not
g43056 not n21538 ; n21538_not
g43057 not n22375 ; n22375_not
g43058 not n26065 ; n26065_not
g43059 not n23671 ; n23671_not
g43060 not n21583 ; n21583_not
g43061 not n22492 ; n22492_not
g43062 not n23554 ; n23554_not
g43063 not n23536 ; n23536_not
g43064 not n26173 ; n26173_not
g43065 not n21592 ; n21592_not
g43066 not n24445 ; n24445_not
g43067 not n23518 ; n23518_not
g43068 not n26164 ; n26164_not
g43069 not n22519 ; n22519_not
g43070 not n24454 ; n24454_not
g43071 not n23509 ; n23509_not
g43072 not n20395 ; n20395_not
g43073 not n23491 ; n23491_not
g43074 not n20386 ; n20386_not
g43075 not n23482 ; n23482_not
g43076 not n22528 ; n22528_not
g43077 not n20359 ; n20359_not
g43078 not n20368 ; n20368_not
g43079 not n22537 ; n22537_not
g43080 not n26218 ; n26218_not
g43081 not n24625 ; n24625_not
g43082 not n24634 ; n24634_not
g43083 not n23608 ; n23608_not
g43084 not n24427 ; n24427_not
g43085 not n22429 ; n22429_not
g43086 not n21565 ; n21565_not
g43087 not n23590 ; n23590_not
g43088 not n26128 ; n26128_not
g43089 not n21574 ; n21574_not
g43090 not n23581 ; n23581_not
g43091 not n22447 ; n22447_not
g43092 not n26137 ; n26137_not
g43093 not n23572 ; n23572_not
g43094 not n20485 ; n20485_not
g43095 not n22456 ; n22456_not
g43096 not n20476 ; n20476_not
g43097 not n26146 ; n26146_not
g43098 not n23563 ; n23563_not
g43099 not n26155 ; n26155_not
g43100 not n20458 ; n20458_not
g43101 not n22474 ; n22474_not
g43102 not n27280 ; n27280_not
g43103 not n22483 ; n22483_not
g43104 not n21862 ; n21862_not
g43105 not n15760 ; n15760_not
g43106 not n11854 ; n11854_not
g43107 not n11638 ; n11638_not
g43108 not n14572 ; n14572_not
g43109 not n14581 ; n14581_not
g43110 not n15751 ; n15751_not
g43111 not n14185 ; n14185_not
g43112 not n11863 ; n11863_not
g43113 not n13096 ; n13096_not
g43114 not n15733 ; n15733_not
g43115 not n18163 ; n18163_not
g43116 not n14590 ; n14590_not
g43117 not n15724 ; n15724_not
g43118 not n15454 ; n15454_not
g43119 not n15715 ; n15715_not
g43120 not n13087 ; n13087_not
g43121 not n18154 ; n18154_not
g43122 not n18082 ; n18082_not
g43123 not n17560 ; n17560_not
g43124 not n13186 ; n13186_not
g43125 not n15841 ; n15841_not
g43126 not n11764 ; n11764_not
g43127 not n11773 ; n11773_not
g43128 not n11782 ; n11782_not
g43129 not n14167 ; n14167_not
g43130 not n15823 ; n15823_not
g43131 not n11467 ; n11467_not
g43132 not n11791 ; n11791_not
g43133 not n13177 ; n13177_not
g43134 not n11809 ; n11809_not
g43135 not n11818 ; n11818_not
g43136 not n18451 ; n18451_not
g43137 not n15814 ; n15814_not
g43138 not n11836 ; n11836_not
g43139 not n18172 ; n18172_not
g43140 not n13168 ; n13168_not
g43141 not n13159 ; n13159_not
g43142 not n11692 ; n11692_not
g43143 not n17632 ; n17632_not
g43144 not n18118 ; n18118_not
g43145 not n15643 ; n15643_not
g43146 not n18109 ; n18109_not
g43147 not n17641 ; n17641_not
g43148 not n11935 ; n11935_not
g43149 not n12619 ; n12619_not
g43150 not n15625 ; n15625_not
g43151 not n17650 ; n17650_not
g43152 not n12880 ; n12880_not
g43153 not n15616 ; n15616_not
g43154 not n11944 ; n11944_not
g43155 not n14635 ; n14635_not
g43156 not n18091 ; n18091_not
g43157 not n14644 ; n14644_not
g43158 not n12925 ; n12925_not
g43159 not n12574 ; n12574_not
g43160 not n11953 ; n11953_not
g43161 not n15580 ; n15580_not
g43162 not n15571 ; n15571_not
g43163 not n18073 ; n18073_not
g43164 not n14653 ; n14653_not
g43165 not n15562 ; n15562_not
g43166 not n16921 ; n16921_not
g43167 not n15706 ; n15706_not
g43168 not n13078 ; n13078_not
g43169 not n13069 ; n13069_not
g43170 not n11881 ; n11881_not
g43171 not n18145 ; n18145_not
g43172 not n11890 ; n11890_not
g43173 not n17605 ; n17605_not
g43174 not n14608 ; n14608_not
g43175 not n18136 ; n18136_not
g43176 not n11908 ; n11908_not
g43177 not n11917 ; n11917_not
g43178 not n14617 ; n14617_not
g43179 not n17614 ; n17614_not
g43180 not n12682 ; n12682_not
g43181 not n15670 ; n15670_not
g43182 not n18127 ; n18127_not
g43183 not n15661 ; n15661_not
g43184 not n17623 ; n17623_not
g43185 not n15652 ; n15652_not
g43186 not n12826 ; n12826_not
g43187 not n13357 ; n13357_not
g43188 not n14491 ; n14491_not
g43189 not n17506 ; n17506_not
g43190 not n13348 ; n13348_not
g43191 not n11476 ; n11476_not
g43192 not n17371 ; n17371_not
g43193 not n17515 ; n17515_not
g43194 not n11287 ; n11287_not
g43195 not n11485 ; n11485_not
g43196 not n14509 ; n14509_not
g43197 not n11494 ; n11494_not
g43198 not n16084 ; n16084_not
g43199 not n13294 ; n13294_not
g43200 not n13285 ; n13285_not
g43201 not n11539 ; n11539_not
g43202 not n11548 ; n11548_not
g43203 not n14518 ; n14518_not
g43204 not n16075 ; n16075_not
g43205 not n14527 ; n14527_not
g43206 not n11557 ; n11557_not
g43207 not n16066 ; n16066_not
g43208 not n16057 ; n16057_not
g43209 not n18244 ; n18244_not
g43210 not n16165 ; n16165_not
g43211 not n11296 ; n11296_not
g43212 not n16156 ; n16156_not
g43213 not n10963 ; n10963_not
g43214 not n14482 ; n14482_not
g43215 not n11359 ; n11359_not
g43216 not n11368 ; n11368_not
g43217 not n16147 ; n16147_not
g43218 not n13375 ; n13375_not
g43219 not n16138 ; n16138_not
g43220 not n18631 ; n18631_not
g43221 not n11377 ; n11377_not
g43222 not n17722 ; n17722_not
g43223 not n16129 ; n16129_not
g43224 not n11386 ; n11386_not
g43225 not n11395 ; n11395_not
g43226 not n11449 ; n11449_not
g43227 not n13366 ; n13366_not
g43228 not n11458 ; n11458_not
g43229 not n18262 ; n18262_not
g43230 not n11656 ; n11656_not
g43231 not n14545 ; n14545_not
g43232 not n11665 ; n11665_not
g43233 not n12844 ; n12844_not
g43234 not n18208 ; n18208_not
g43235 not n11674 ; n11674_not
g43236 not n15922 ; n15922_not
g43237 not n11683 ; n11683_not
g43238 not n15913 ; n15913_not
g43239 not n15904 ; n15904_not
g43240 not n17551 ; n17551_not
g43241 not n11719 ; n11719_not
g43242 not n11728 ; n11728_not
g43243 not n11746 ; n11746_not
g43244 not n14554 ; n14554_not
g43245 not n15850 ; n15850_not
g43246 not n14563 ; n14563_not
g43247 not n15832 ; n15832_not
g43248 not n16039 ; n16039_not
g43249 not n11566 ; n11566_not
g43250 not n13276 ; n13276_not
g43251 not n13267 ; n13267_not
g43252 not n18622 ; n18622_not
g43253 not n11575 ; n11575_not
g43254 not n18613 ; n18613_not
g43255 not n11584 ; n11584_not
g43256 not n17533 ; n17533_not
g43257 not n14536 ; n14536_not
g43258 not n11593 ; n11593_not
g43259 not n18226 ; n18226_not
g43260 not n13258 ; n13258_not
g43261 not n15940 ; n15940_not
g43262 not n11629 ; n11629_not
g43263 not n11647 ; n11647_not
g43264 not n13249 ; n13249_not
g43265 not n15931 ; n15931_not
g43266 not n14824 ; n14824_not
g43267 not n15238 ; n15238_not
g43268 not n15193 ; n15193_not
g43269 not n12493 ; n12493_not
g43270 not n12484 ; n12484_not
g43271 not n12772 ; n12772_not
g43272 not n14833 ; n14833_not
g43273 not n15184 ; n15184_not
g43274 not n15175 ; n15175_not
g43275 not n14842 ; n14842_not
g43276 not n12529 ; n12529_not
g43277 not n12277 ; n12277_not
g43278 not n12538 ; n12538_not
g43279 not n15166 ; n15166_not
g43280 not n14851 ; n14851_not
g43281 not n12547 ; n12547_not
g43282 not n12763 ; n12763_not
g43283 not n12556 ; n12556_not
g43284 not n15148 ; n15148_not
g43285 not n15139 ; n15139_not
g43286 not n12439 ; n12439_not
g43287 not n12448 ; n12448_not
g43288 not n14941 ; n14941_not
g43289 not n18514 ; n18514_not
g43290 not n14806 ; n14806_not
g43291 not n17821 ; n17821_not
g43292 not n12808 ; n12808_not
g43293 not n15283 ; n15283_not
g43294 not n12457 ; n12457_not
g43295 not n14680 ; n14680_not
g43296 not n17830 ; n17830_not
g43297 not n14815 ; n14815_not
g43298 not n15274 ; n15274_not
g43299 not n15265 ; n15265_not
g43300 not n12466 ; n12466_not
g43301 not n12790 ; n12790_not
g43302 not n15256 ; n15256_not
g43303 not n15247 ; n15247_not
g43304 not n12475 ; n12475_not
g43305 not n12637 ; n12637_not
g43306 not n12646 ; n12646_not
g43307 not n12736 ; n12736_not
g43308 not n12655 ; n12655_not
g43309 not n14950 ; n14950_not
g43310 not n17920 ; n17920_not
g43311 not n17902 ; n17902_not
g43312 not n14905 ; n14905_not
g43313 not n12727 ; n12727_not
g43314 not n12664 ; n12664_not
g43315 not n14932 ; n14932_not
g43316 not n12673 ; n12673_not
g43317 not n14923 ; n14923_not
g43318 not n12718 ; n12718_not
g43319 not n12709 ; n12709_not
g43320 not n12394 ; n12394_not
g43321 not n12691 ; n12691_not
g43322 not n14275 ; n14275_not
g43323 not n14752 ; n14752_not
g43324 not n12565 ; n12565_not
g43325 not n15094 ; n15094_not
g43326 not n14365 ; n14365_not
g43327 not n14860 ; n14860_not
g43328 not n15085 ; n15085_not
g43329 not n12754 ; n12754_not
g43330 not n15076 ; n15076_not
g43331 not n12592 ; n12592_not
g43332 not n15067 ; n15067_not
g43333 not n15058 ; n15058_not
g43334 not n15049 ; n15049_not
g43335 not n12628 ; n12628_not
g43336 not n14707 ; n14707_not
g43337 not n11926 ; n11926_not
g43338 not n12376 ; n12376_not
g43339 not n12745 ; n12745_not
g43340 not n17317 ; n17317_not
g43341 not n12943 ; n12943_not
g43342 not n12952 ; n12952_not
g43343 not n17731 ; n17731_not
g43344 not n18037 ; n18037_not
g43345 not n18028 ; n18028_not
g43346 not n15490 ; n15490_not
g43347 not n15481 ; n15481_not
g43348 not n14716 ; n14716_not
g43349 not n12934 ; n12934_not
g43350 not n12079 ; n12079_not
g43351 not n17470 ; n17470_not
g43352 not n15472 ; n15472_not
g43353 not n14725 ; n14725_not
g43354 not n12916 ; n12916_not
g43355 not n12907 ; n12907_not
g43356 not n11827 ; n11827_not
g43357 not n15463 ; n15463_not
g43358 not n12169 ; n12169_not
g43359 not n11962 ; n11962_not
g43360 not n15517 ; n15517_not
g43361 not n14662 ; n14662_not
g43362 not n18550 ; n18550_not
g43363 not n15553 ; n15553_not
g43364 not n18064 ; n18064_not
g43365 not n15544 ; n15544_not
g43366 not n11980 ; n11980_not
g43367 not n15535 ; n15535_not
g43368 not n14428 ; n14428_not
g43369 not n17704 ; n17704_not
g43370 not n12970 ; n12970_not
g43371 not n15526 ; n15526_not
g43372 not n18046 ; n18046_not
g43373 not n17713 ; n17713_not
g43374 not n15508 ; n15508_not
g43375 not n15382 ; n15382_not
g43376 not n12367 ; n12367_not
g43377 not n12358 ; n12358_not
g43378 not n15373 ; n15373_not
g43379 not n12835 ; n12835_not
g43380 not n15364 ; n15364_not
g43381 not n12385 ; n12385_not
g43382 not n15355 ; n15355_not
g43383 not n15346 ; n15346_not
g43384 not n15337 ; n15337_not
g43385 not n12817 ; n12817_not
g43386 not n15328 ; n15328_not
g43387 not n15319 ; n15319_not
g43388 not n18523 ; n18523_not
g43389 not n17812 ; n17812_not
g43390 not n12178 ; n12178_not
g43391 not n12187 ; n12187_not
g43392 not n14257 ; n14257_not
g43393 not n14734 ; n14734_not
g43394 not n15445 ; n15445_not
g43395 not n15436 ; n15436_not
g43396 not n14743 ; n14743_not
g43397 not n15418 ; n15418_not
g43398 not n12259 ; n12259_not
g43399 not n12268 ; n12268_not
g43400 not n12286 ; n12286_not
g43401 not n12871 ; n12871_not
g43402 not n14761 ; n14761_not
g43403 not n15391 ; n15391_not
g43404 not n12862 ; n12862_not
g43405 not n12295 ; n12295_not
g43406 not n14770 ; n14770_not
g43407 not n12349 ; n12349_not
g43408 not n10648 ; n10648_not
g43409 not n17245 ; n17245_not
g43410 not n14248 ; n14248_not
g43411 not n10657 ; n10657_not
g43412 not n14239 ; n14239_not
g43413 not n13672 ; n13672_not
g43414 not n10666 ; n10666_not
g43415 not n13663 ; n13663_not
g43416 not n13924 ; n13924_not
g43417 not n16633 ; n16633_not
g43418 not n10675 ; n10675_not
g43419 not n16381 ; n16381_not
g43420 not n13654 ; n13654_not
g43421 not n14266 ; n14266_not
g43422 not n16624 ; n16624_not
g43423 not n17263 ; n17263_not
g43424 not n13645 ; n13645_not
g43425 not n13447 ; n13447_not
g43426 not n16606 ; n16606_not
g43427 not n17236 ; n17236_not
g43428 not n13735 ; n13735_not
g43429 not n18433 ; n18433_not
g43430 not n16714 ; n16714_not
g43431 not n10576 ; n10576_not
g43432 not n14176 ; n14176_not
g43433 not n13717 ; n13717_not
g43434 not n13708 ; n13708_not
g43435 not n18424 ; n18424_not
g43436 not n17209 ; n17209_not
g43437 not n10594 ; n10594_not
g43438 not n17218 ; n17218_not
g43439 not n13690 ; n13690_not
g43440 not n18415 ; n18415_not
g43441 not n18406 ; n18406_not
g43442 not n14194 ; n14194_not
g43443 not n13681 ; n13681_not
g43444 not n16651 ; n16651_not
g43445 not n16642 ; n16642_not
g43446 not n10639 ; n10639_not
g43447 not n13582 ; n13582_not
g43448 not n18370 ; n18370_not
g43449 not n16543 ; n16543_not
g43450 not n16534 ; n16534_not
g43451 not n14293 ; n14293_not
g43452 not n17344 ; n17344_not
g43453 not n13573 ; n13573_not
g43454 not n18361 ; n18361_not
g43455 not n10783 ; n10783_not
g43456 not n14329 ; n14329_not
g43457 not n16525 ; n16525_not
g43458 not n10819 ; n10819_not
g43459 not n16516 ; n16516_not
g43460 not n17353 ; n17353_not
g43461 not n14338 ; n14338_not
g43462 not n16507 ; n16507_not
g43463 not n10837 ; n10837_not
g43464 not n10828 ; n10828_not
g43465 not n14347 ; n14347_not
g43466 not n10792 ; n10792_not
g43467 not n10846 ; n10846_not
g43468 not n13564 ; n13564_not
g43469 not n10693 ; n10693_not
g43470 not n17272 ; n17272_not
g43471 not n13618 ; n13618_not
g43472 not n17281 ; n17281_not
g43473 not n13627 ; n13627_not
g43474 not n10738 ; n10738_not
g43475 not n10558 ; n10558_not
g43476 not n13609 ; n13609_not
g43477 not n10747 ; n10747_not
g43478 not n17290 ; n17290_not
g43479 not n16570 ; n16570_not
g43480 not n13591 ; n13591_not
g43481 not n14284 ; n14284_not
g43482 not n16552 ; n16552_not
g43483 not n10765 ; n10765_not
g43484 not n17326 ; n17326_not
g43485 not n10774 ; n10774_not
g43486 not n17047 ; n17047_not
g43487 not n13816 ; n13816_not
g43488 not n13807 ; n13807_not
g43489 not n16831 ; n16831_not
g43490 not n13951 ; n13951_not
g43491 not n17065 ; n17065_not
g43492 not n17056 ; n17056_not
g43493 not n16813 ; n16813_not
g43494 not n16561 ; n16561_not
g43495 not n17074 ; n17074_not
g43496 not n16804 ; n16804_not
g43497 not n17083 ; n17083_not
g43498 not n14077 ; n14077_not
g43499 not n13780 ; n13780_not
g43500 not n17092 ; n17092_not
g43501 not n10099 ; n10099_not
g43502 not n10189 ; n10189_not
g43503 not n10198 ; n10198_not
g43504 not n10279 ; n10279_not
g43505 not n13915 ; n13915_not
g43506 not n13906 ; n13906_not
g43507 not n13870 ; n13870_not
g43508 not n16930 ; n16930_not
g43509 not n16912 ; n16912_not
g43510 not n16840 ; n16840_not
g43511 not n13933 ; n13933_not
g43512 not n13852 ; n13852_not
g43513 not n16903 ; n16903_not
g43514 not n13843 ; n13843_not
g43515 not n13834 ; n13834_not
g43516 not n16723 ; n16723_not
g43517 not n13474 ; n13474_not
g43518 not n17029 ; n17029_not
g43519 not n17038 ; n17038_not
g43520 not n13960 ; n13960_not
g43521 not n17146 ; n17146_not
g43522 not n10495 ; n10495_not
g43523 not n16750 ; n16750_not
g43524 not n14149 ; n14149_not
g43525 not n14158 ; n14158_not
g43526 not n16741 ; n16741_not
g43527 not n13753 ; n13753_not
g43528 not n17173 ; n17173_not
g43529 not n13744 ; n13744_not
g43530 not n17164 ; n17164_not
g43531 not n16426 ; n16426_not
g43532 not n16732 ; n16732_not
g43533 not n10549 ; n10549_not
g43534 not n17182 ; n17182_not
g43535 not n16615 ; n16615_not
g43536 not n10567 ; n10567_not
g43537 not n17191 ; n17191_not
g43538 not n10288 ; n10288_not
g43539 not n14086 ; n14086_not
g43540 not n10297 ; n10297_not
g43541 not n17119 ; n17119_not
g43542 not n14095 ; n14095_not
g43543 not n10369 ; n10369_not
g43544 not n10378 ; n10378_not
g43545 not n10387 ; n10387_not
g43546 not n17128 ; n17128_not
g43547 not n17137 ; n17137_not
g43548 not n13762 ; n13762_not
g43549 not n10459 ; n10459_not
g43550 not n10468 ; n10468_not
g43551 not n10477 ; n10477_not
g43552 not n17155 ; n17155_not
g43553 not n10486 ; n10486_not
g43554 not n14455 ; n14455_not
g43555 not n14383 ; n14383_not
g43556 not n17407 ; n17407_not
g43557 not n10927 ; n10927_not
g43558 not n14419 ; n14419_not
g43559 not n16417 ; n16417_not
g43560 not n13519 ; n13519_not
g43561 not n16246 ; n16246_not
g43562 not n16462 ; n16462_not
g43563 not n17452 ; n17452_not
g43564 not n18334 ; n18334_not
g43565 not n13528 ; n13528_not
g43566 not n16237 ; n16237_not
g43567 not n10873 ; n10873_not
g43568 not n10981 ; n10981_not
g43569 not n11179 ; n11179_not
g43570 not n16471 ; n16471_not
g43571 not n16309 ; n16309_not
g43572 not n10864 ; n10864_not
g43573 not n18280 ; n18280_not
g43574 not n14437 ; n14437_not
g43575 not n14464 ; n14464_not
g43576 not n14473 ; n14473_not
g43577 not n11188 ; n11188_not
g43578 not n13438 ; n13438_not
g43579 not n14392 ; n14392_not
g43580 not n10990 ; n10990_not
g43581 not n13429 ; n13429_not
g43582 not n17434 ; n17434_not
g43583 not n13483 ; n13483_not
g43584 not n16273 ; n16273_not
g43585 not n16444 ; n16444_not
g43586 not n16453 ; n16453_not
g43587 not n18325 ; n18325_not
g43588 not n16435 ; n16435_not
g43589 not n13492 ; n13492_not
g43590 not n16264 ; n16264_not
g43591 not n10891 ; n10891_not
g43592 not n17416 ; n17416_not
g43593 not n10729 ; n10729_not
g43594 not n10909 ; n10909_not
g43595 not n11098 ; n11098_not
g43596 not n16282 ; n16282_not
g43597 not n10882 ; n10882_not
g43598 not n16291 ; n16291_not
g43599 not n13456 ; n13456_not
g43600 not n18307 ; n18307_not
g43601 not n11269 ; n11269_not
g43602 not n11278 ; n11278_not
g43603 not n16480 ; n16480_not
g43604 not n16174 ; n16174_not
g43605 not n10855 ; n10855_not
g43606 not n17461 ; n17461_not
g43607 not n16183 ; n16183_not
g43608 not n10918 ; n10918_not
g43609 not n13555 ; n13555_not
g43610 not n10945 ; n10945_not
g43611 not n13384 ; n13384_not
g43612 not n16372 ; n16372_not
g43613 not n14356 ; n14356_not
g43614 not n14446 ; n14446_not
g43615 not n16363 ; n16363_not
g43616 not n10954 ; n10954_not
g43617 not n18352 ; n18352_not
g43618 not n17362 ; n17362_not
g43619 not n13393 ; n13393_not
g43620 not n10972 ; n10972_not
g43621 not n18343 ; n18343_not
g43622 not n16219 ; n16219_not
g43623 not n11197 ; n11197_not
g43624 not n10756 ; n10756_not
g43625 not n16228 ; n16228_not
g43626 not n14374 ; n14374_not
g43627 not n16327 ; n16327_not
g43628 not n13546 ; n13546_not
g43629 not n16345 ; n16345_not
g43630 not n10936 ; n10936_not
g43631 not n17380 ; n17380_not
g43632 not n16390 ; n16390_not
g43633 not n18019 ; n18019_not
g43634 not n17633 ; n17633_not
g43635 not n23375 ; n23375_not
g43636 not n23366 ; n23366_not
g43637 not n18236 ; n18236_not
g43638 not n23852 ; n23852_not
g43639 not n14096 ; n14096_not
g43640 not n13844 ; n13844_not
g43641 not n23681 ; n23681_not
g43642 not n14519 ; n14519_not
g43643 not n14825 ; n14825_not
g43644 not n13673 ; n13673_not
g43645 not n23348 ; n23348_not
g43646 not n18227 ; n18227_not
g43647 not n14447 ; n14447_not
g43648 not n14456 ; n14456_not
g43649 not n14816 ; n14816_not
g43650 not n23555 ; n23555_not
g43651 not n14528 ; n14528_not
g43652 not n18290 ; n18290_not
g43653 not n14807 ; n14807_not
g43654 not n23780 ; n23780_not
g43655 not n18245 ; n18245_not
g43656 not n20369 ; n20369_not
g43657 not n23276 ; n23276_not
g43658 not n13943 ; n13943_not
g43659 not n14474 ; n14474_not
g43660 not n17930 ; n17930_not
g43661 not n23294 ; n23294_not
g43662 not n13529 ; n13529_not
g43663 not n13952 ; n13952_not
g43664 not n23285 ; n23285_not
g43665 not n14384 ; n14384_not
g43666 not n14870 ; n14870_not
g43667 not n18263 ; n18263_not
g43668 not n13961 ; n13961_not
g43669 not n14492 ; n14492_not
g43670 not n18281 ; n18281_not
g43671 not n14861 ; n14861_not
g43672 not n20396 ; n20396_not
g43673 not n13547 ; n13547_not
g43674 not n24185 ; n24185_not
g43675 not n17921 ; n17921_not
g43676 not n24176 ; n24176_not
g43677 not n13907 ; n13907_not
g43678 not n13916 ; n13916_not
g43679 not n18272 ; n18272_not
g43680 not n23726 ; n23726_not
g43681 not n23483 ; n23483_not
g43682 not n24158 ; n24158_not
g43683 not n14483 ; n14483_not
g43684 not n23735 ; n23735_not
g43685 not n23744 ; n23744_not
g43686 not n13934 ; n13934_not
g43687 not n13925 ; n13925_not
g43688 not n23708 ; n23708_not
g43689 not n23645 ; n23645_not
g43690 not n14078 ; n14078_not
g43691 not n23339 ; n23339_not
g43692 not n14843 ; n14843_not
g43693 not n23771 ; n23771_not
g43694 not n20387 ; n20387_not
g43695 not n13655 ; n13655_not
g43696 not n14348 ; n14348_not
g43697 not n14834 ; n14834_not
g43698 not n24068 ; n24068_not
g43699 not n20378 ; n20378_not
g43700 not n23357 ; n23357_not
g43701 not n18254 ; n18254_not
g43702 not n13970 ; n13970_not
g43703 not n13556 ; n13556_not
g43704 not n23717 ; n23717_not
g43705 not n14852 ; n14852_not
g43706 not n18065 ; n18065_not
g43707 not n24095 ; n24095_not
g43708 not n24086 ; n24086_not
g43709 not n13592 ; n13592_not
g43710 not n23609 ; n23609_not
g43711 not n13637 ; n13637_not
g43712 not n14069 ; n14069_not
g43713 not n23762 ; n23762_not
g43714 not n24077 ; n24077_not
g43715 not n14645 ; n14645_not
g43716 not n14375 ; n14375_not
g43717 not n23825 ; n23825_not
g43718 not n23843 ; n23843_not
g43719 not n23942 ; n23942_not
g43720 not n18092 ; n18092_not
g43721 not n14636 ; n14636_not
g43722 not n14573 ; n14573_not
g43723 not n23564 ; n23564_not
g43724 not n23573 ; n23573_not
g43725 not n18083 ; n18083_not
g43726 not n20288 ; n20288_not
g43727 not n14276 ; n14276_not
g43728 not n17912 ; n17912_not
g43729 not n14672 ; n14672_not
g43730 not n23519 ; n23519_not
g43731 not n23528 ; n23528_not
g43732 not n14663 ; n14663_not
g43733 not n23960 ; n23960_not
g43734 not n18173 ; n18173_not
g43735 not n14465 ; n14465_not
g43736 not n23834 ; n23834_not
g43737 not n23951 ; n23951_not
g43738 not n18074 ; n18074_not
g43739 not n14654 ; n14654_not
g43740 not n23537 ; n23537_not
g43741 not n23546 ; n23546_not
g43742 not n14366 ; n14366_not
g43743 not n18164 ; n18164_not
g43744 not n18137 ; n18137_not
g43745 not n23861 ; n23861_not
g43746 not n14609 ; n14609_not
g43747 not n17831 ; n17831_not
g43748 not n23591 ; n23591_not
g43749 not n14339 ; n14339_not
g43750 not n18146 ; n18146_not
g43751 not n18155 ; n18155_not
g43752 not n23384 ; n23384_not
g43753 not n18353 ; n18353_not
g43754 not n14285 ; n14285_not
g43755 not n23627 ; n23627_not
g43756 not n23618 ; n23618_not
g43757 not n18344 ; n18344_not
g43758 not n18119 ; n18119_not
g43759 not n23924 ; n23924_not
g43760 not n14582 ; n14582_not
g43761 not n18362 ; n18362_not
g43762 not n14618 ; n14618_not
g43763 not n23906 ; n23906_not
g43764 not n18128 ; n18128_not
g43765 not n14762 ; n14762_not
g43766 not n23672 ; n23672_not
g43767 not n14177 ; n14177_not
g43768 not n13808 ; n13808_not
g43769 not n23438 ; n23438_not
g43770 not n18308 ; n18308_not
g43771 not n14753 ; n14753_not
g43772 not n18425 ; n18425_not
g43773 not n23663 ; n23663_not
g43774 not n14744 ; n14744_not
g43775 not n14735 ; n14735_not
g43776 not n14186 ; n14186_not
g43777 not n14195 ; n14195_not
g43778 not n14546 ; n14546_not
g43779 not n23465 ; n23465_not
g43780 not n14537 ; n14537_not
g43781 not n18434 ; n18434_not
g43782 not n14438 ; n14438_not
g43783 not n14159 ; n14159_not
g43784 not n23393 ; n23393_not
g43785 not n14780 ; n14780_not
g43786 not n14771 ; n14771_not
g43787 not n18209 ; n18209_not
g43788 not n23429 ; n23429_not
g43789 not n14168 ; n14168_not
g43790 not n14393 ; n14393_not
g43791 not n18326 ; n18326_not
g43792 not n18038 ; n18038_not
g43793 not n14564 ; n14564_not
g43794 not n18047 ; n18047_not
g43795 not n18182 ; n18182_not
g43796 not n23492 ; n23492_not
g43797 not n20297 ; n20297_not
g43798 not n14267 ; n14267_not
g43799 not n14690 ; n14690_not
g43800 not n23636 ; n23636_not
g43801 not n14258 ; n14258_not
g43802 not n14726 ; n14726_not
g43803 not n18407 ; n18407_not
g43804 not n18191 ; n18191_not
g43805 not n23474 ; n23474_not
g43806 not n23654 ; n23654_not
g43807 not n14717 ; n14717_not
g43808 not n19910 ; n19910_not
g43809 not n14555 ; n14555_not
g43810 not n14708 ; n14708_not
g43811 not n14249 ; n14249_not
g43812 not n20198 ; n20198_not
g43813 not n18029 ; n18029_not
g43814 not n21935 ; n21935_not
g43815 not n21944 ; n21944_not
g43816 not n16463 ; n16463_not
g43817 not n21953 ; n21953_not
g43818 not n17408 ; n17408_not
g43819 not n16454 ; n16454_not
g43820 not n21971 ; n21971_not
g43821 not n17417 ; n17417_not
g43822 not n17426 ; n17426_not
g43823 not n21746 ; n21746_not
g43824 not n16445 ; n16445_not
g43825 not n17435 ; n17435_not
g43826 not n16436 ; n16436_not
g43827 not n16418 ; n16418_not
g43828 not n17453 ; n17453_not
g43829 not n17093 ; n17093_not
g43830 not n16409 ; n16409_not
g43831 not n21764 ; n21764_not
g43832 not n16391 ; n16391_not
g43833 not n21782 ; n21782_not
g43834 not n16382 ; n16382_not
g43835 not n15932 ; n15932_not
g43836 not n16364 ; n16364_not
g43837 not n21980 ; n21980_not
g43838 not n20990 ; n20990_not
g43839 not n16346 ; n16346_not
g43840 not n16337 ; n16337_not
g43841 not n16328 ; n16328_not
g43842 not n15905 ; n15905_not
g43843 not n21845 ; n21845_not
g43844 not n21089 ; n21089_not
g43845 not n17336 ; n17336_not
g43846 not n17345 ; n17345_not
g43847 not n20873 ; n20873_not
g43848 not n16526 ; n16526_not
g43849 not n17354 ; n17354_not
g43850 not n16508 ; n16508_not
g43851 not n21863 ; n21863_not
g43852 not n17363 ; n17363_not
g43853 not n21881 ; n21881_not
g43854 not n21890 ; n21890_not
g43855 not n16490 ; n16490_not
g43856 not n21692 ; n21692_not
g43857 not n21908 ; n21908_not
g43858 not n17372 ; n17372_not
g43859 not n16481 ; n16481_not
g43860 not n17381 ; n17381_not
g43861 not n21917 ; n21917_not
g43862 not n17048 ; n17048_not
g43863 not n17390 ; n17390_not
g43864 not n16472 ; n16472_not
g43865 not n16292 ; n16292_not
g43866 not n20927 ; n20927_not
g43867 not n15419 ; n15419_not
g43868 not n22169 ; n22169_not
g43869 not n21926 ; n21926_not
g43870 not n20918 ; n20918_not
g43871 not n22178 ; n22178_not
g43872 not n17507 ; n17507_not
g43873 not n16094 ; n16094_not
g43874 not n22187 ; n22187_not
g43875 not n20909 ; n20909_not
g43876 not n16085 ; n16085_not
g43877 not n17525 ; n17525_not
g43878 not n22196 ; n22196_not
g43879 not n16076 ; n16076_not
g43880 not n16067 ; n16067_not
g43881 not n16058 ; n16058_not
g43882 not n20891 ; n20891_not
g43883 not n16049 ; n16049_not
g43884 not n22097 ; n22097_not
g43885 not n22259 ; n22259_not
g43886 not n22268 ; n22268_not
g43887 not n15950 ; n15950_not
g43888 not n20882 ; n20882_not
g43889 not n17534 ; n17534_not
g43890 not n22286 ; n22286_not
g43891 not n22088 ; n22088_not
g43892 not n16283 ; n16283_not
g43893 not n20972 ; n20972_not
g43894 not n16274 ; n16274_not
g43895 not n20738 ; n20738_not
g43896 not n16265 ; n16265_not
g43897 not n20963 ; n20963_not
g43898 not n17471 ; n17471_not
g43899 not n16256 ; n16256_not
g43900 not n16247 ; n16247_not
g43901 not n20954 ; n20954_not
g43902 not n16238 ; n16238_not
g43903 not n16229 ; n16229_not
g43904 not n17480 ; n17480_not
g43905 not n20945 ; n20945_not
g43906 not n16184 ; n16184_not
g43907 not n16175 ; n16175_not
g43908 not n20936 ; n20936_not
g43909 not n16166 ; n16166_not
g43910 not n16157 ; n16157_not
g43911 not n16148 ; n16148_not
g43912 not n16139 ; n16139_not
g43913 not n21278 ; n21278_not
g43914 not n16814 ; n16814_not
g43915 not n17075 ; n17075_not
g43916 not n21269 ; n21269_not
g43917 not n16805 ; n16805_not
g43918 not n21539 ; n21539_not
g43919 not n17084 ; n17084_not
g43920 not n21485 ; n21485_not
g43921 not n21548 ; n21548_not
g43922 not n21557 ; n21557_not
g43923 not n21566 ; n21566_not
g43924 not n16760 ; n16760_not
g43925 not n21584 ; n21584_not
g43926 not n17129 ; n17129_not
g43927 not n17138 ; n17138_not
g43928 not n21593 ; n21593_not
g43929 not n17147 ; n17147_not
g43930 not n17156 ; n17156_not
g43931 not n16751 ; n16751_not
g43932 not n16742 ; n16742_not
g43933 not n17165 ; n17165_not
g43934 not n17174 ; n17174_not
g43935 not n16733 ; n16733_not
g43936 not n17183 ; n17183_not
g43937 not n21629 ; n21629_not
g43938 not n16940 ; n16940_not
g43939 not n21359 ; n21359_not
g43940 not n16931 ; n16931_not
g43941 not n21377 ; n21377_not
g43942 not n16922 ; n16922_not
g43943 not n16913 ; n16913_not
g43944 not n21395 ; n21395_not
g43945 not n16904 ; n16904_not
g43946 not n21449 ; n21449_not
g43947 not n21467 ; n21467_not
g43948 not n16850 ; n16850_not
g43949 not n21476 ; n21476_not
g43950 not n16841 ; n16841_not
g43951 not n16706 ; n16706_not
g43952 not n16652 ; n16652_not
g43953 not n16832 ; n16832_not
g43954 not n17039 ; n17039_not
g43955 not n21494 ; n21494_not
g43956 not n21287 ; n21287_not
g43957 not n17057 ; n17057_not
g43958 not n17066 ; n17066_not
g43959 not n16823 ; n16823_not
g43960 not n21728 ; n21728_not
g43961 not n16625 ; n16625_not
g43962 not n21737 ; n21737_not
g43963 not n17264 ; n17264_not
g43964 not n16607 ; n16607_not
g43965 not n21755 ; n21755_not
g43966 not n16580 ; n16580_not
g43967 not n17282 ; n17282_not
g43968 not n17228 ; n17228_not
g43969 not n21791 ; n21791_not
g43970 not n16571 ; n16571_not
g43971 not n17291 ; n17291_not
g43972 not n16562 ; n16562_not
g43973 not n21809 ; n21809_not
g43974 not n16553 ; n16553_not
g43975 not n17309 ; n17309_not
g43976 not n17318 ; n17318_not
g43977 not n16544 ; n16544_not
g43978 not n17327 ; n17327_not
g43979 not n21827 ; n21827_not
g43980 not n21098 ; n21098_not
g43981 not n21458 ; n21458_not
g43982 not n17192 ; n17192_not
g43983 not n16715 ; n16715_not
g43984 not n16616 ; n16616_not
g43985 not n21638 ; n21638_not
g43986 not n21647 ; n21647_not
g43987 not n21197 ; n21197_not
g43988 not n21656 ; n21656_not
g43989 not n16670 ; n16670_not
g43990 not n21674 ; n21674_not
g43991 not n21188 ; n21188_not
g43992 not n17219 ; n17219_not
g43993 not n21179 ; n21179_not
g43994 not n16661 ; n16661_not
g43995 not n17237 ; n17237_not
g43996 not n21719 ; n21719_not
g43997 not n17246 ; n17246_not
g43998 not n16643 ; n16643_not
g43999 not n16634 ; n16634_not
g44000 not n15284 ; n15284_not
g44001 not n20576 ; n20576_not
g44002 not n22907 ; n22907_not
g44003 not n22673 ; n22673_not
g44004 not n20567 ; n20567_not
g44005 not n22916 ; n22916_not
g44006 not n15392 ; n15392_not
g44007 not n22925 ; n22925_not
g44008 not n22934 ; n22934_not
g44009 not n15383 ; n15383_not
g44010 not n22952 ; n22952_not
g44011 not n22961 ; n22961_not
g44012 not n20549 ; n20549_not
g44013 not n22808 ; n22808_not
g44014 not n22970 ; n22970_not
g44015 not n15347 ; n15347_not
g44016 not n15365 ; n15365_not
g44017 not n22754 ; n22754_not
g44018 not n15356 ; n15356_not
g44019 not n15338 ; n15338_not
g44020 not n15329 ; n15329_not
g44021 not n22781 ; n22781_not
g44022 not n15527 ; n15527_not
g44023 not n17705 ; n17705_not
g44024 not n15518 ; n15518_not
g44025 not n15509 ; n15509_not
g44026 not n17723 ; n17723_not
g44027 not n15491 ; n15491_not
g44028 not n17732 ; n17732_not
g44029 not n22727 ; n22727_not
g44030 not n15482 ; n15482_not
g44031 not n15239 ; n15239_not
g44032 not n22817 ; n22817_not
g44033 not n22826 ; n22826_not
g44034 not n17750 ; n17750_not
g44035 not n22583 ; n22583_not
g44036 not n22835 ; n22835_not
g44037 not n15464 ; n15464_not
g44038 not n22844 ; n22844_not
g44039 not n15455 ; n15455_not
g44040 not n20594 ; n20594_not
g44041 not n22853 ; n22853_not
g44042 not n22871 ; n22871_not
g44043 not n20585 ; n20585_not
g44044 not n15446 ; n15446_not
g44045 not n15086 ; n15086_not
g44046 not n15077 ; n15077_not
g44047 not n20459 ; n20459_not
g44048 not n15068 ; n15068_not
g44049 not n23159 ; n23159_not
g44050 not n23168 ; n23168_not
g44051 not n23177 ; n23177_not
g44052 not n23186 ; n23186_not
g44053 not n23195 ; n23195_not
g44054 not n14960 ; n14960_not
g44055 not n14951 ; n14951_not
g44056 not n14942 ; n14942_not
g44057 not n17903 ; n17903_not
g44058 not n14924 ; n14924_not
g44059 not n14933 ; n14933_not
g44060 not n23258 ; n23258_not
g44061 not n23249 ; n23249_not
g44062 not n14915 ; n14915_not
g44063 not n14681 ; n14681_not
g44064 not n23267 ; n23267_not
g44065 not n14906 ; n14906_not
g44066 not n17813 ; n17813_not
g44067 not n15293 ; n15293_not
g44068 not n15275 ; n15275_not
g44069 not n15266 ; n15266_not
g44070 not n15257 ; n15257_not
g44071 not n23069 ; n23069_not
g44072 not n15248 ; n15248_not
g44073 not n23078 ; n23078_not
g44074 not n17840 ; n17840_not
g44075 not n15194 ; n15194_not
g44076 not n20495 ; n20495_not
g44077 not n23096 ; n23096_not
g44078 not n23087 ; n23087_not
g44079 not n15185 ; n15185_not
g44080 not n15176 ; n15176_not
g44081 not n22943 ; n22943_not
g44082 not n15167 ; n15167_not
g44083 not n15158 ; n15158_not
g44084 not n20477 ; n20477_not
g44085 not n15149 ; n15149_not
g44086 not n15095 ; n15095_not
g44087 not n17570 ; n17570_not
g44088 not n15815 ; n15815_not
g44089 not n15770 ; n15770_not
g44090 not n22448 ; n22448_not
g44091 not n22457 ; n22457_not
g44092 not n22466 ; n22466_not
g44093 not n15761 ; n15761_not
g44094 not n22475 ; n22475_not
g44095 not n22484 ; n22484_not
g44096 not n15752 ; n15752_not
g44097 not n15743 ; n15743_not
g44098 not n20783 ; n20783_not
g44099 not n15734 ; n15734_not
g44100 not n17273 ; n17273_not
g44101 not n15725 ; n15725_not
g44102 not n15716 ; n15716_not
g44103 not n20774 ; n20774_not
g44104 not n22529 ; n22529_not
g44105 not n22538 ; n22538_not
g44106 not n20765 ; n20765_not
g44107 not n15707 ; n15707_not
g44108 not n22547 ; n22547_not
g44109 not n22556 ; n22556_not
g44110 not n15941 ; n15941_not
g44111 not n22295 ; n22295_not
g44112 not n15914 ; n15914_not
g44113 not n17543 ; n17543_not
g44114 not n22277 ; n22277_not
g44115 not n15923 ; n15923_not
g44116 not n20855 ; n20855_not
g44117 not n15536 ; n15536_not
g44118 not n22358 ; n22358_not
g44119 not n15608 ; n15608_not
g44120 not n22367 ; n22367_not
g44121 not n17552 ; n17552_not
g44122 not n15860 ; n15860_not
g44123 not n22376 ; n22376_not
g44124 not n22385 ; n22385_not
g44125 not n20837 ; n20837_not
g44126 not n22394 ; n22394_not
g44127 not n20828 ; n20828_not
g44128 not n15842 ; n15842_not
g44129 not n17561 ; n17561_not
g44130 not n15833 ; n15833_not
g44131 not n20819 ; n20819_not
g44132 not n15824 ; n15824_not
g44133 not n22655 ; n22655_not
g44134 not n15590 ; n15590_not
g44135 not n17660 ; n17660_not
g44136 not n22664 ; n22664_not
g44137 not n15581 ; n15581_not
g44138 not n20693 ; n20693_not
g44139 not n22682 ; n22682_not
g44140 not n22691 ; n22691_not
g44141 not n22646 ; n22646_not
g44142 not n20684 ; n20684_not
g44143 not n15572 ; n15572_not
g44144 not n22637 ; n22637_not
g44145 not n22718 ; n22718_not
g44146 not n15563 ; n15563_not
g44147 not n20675 ; n20675_not
g44148 not n22736 ; n22736_not
g44149 not n15554 ; n15554_not
g44150 not n20666 ; n20666_not
g44151 not n15545 ; n15545_not
g44152 not n20648 ; n20648_not
g44153 not n22772 ; n22772_not
g44154 not n20756 ; n20756_not
g44155 not n20639 ; n20639_not
g44156 not n22565 ; n22565_not
g44157 not n22574 ; n22574_not
g44158 not n17606 ; n17606_not
g44159 not n22592 ; n22592_not
g44160 not n20747 ; n20747_not
g44161 not n17255 ; n17255_not
g44162 not n17615 ; n17615_not
g44163 not n15653 ; n15653_not
g44164 not n15662 ; n15662_not
g44165 not n17624 ; n17624_not
g44166 not n20729 ; n20729_not
g44167 not n22619 ; n22619_not
g44168 not n22628 ; n22628_not
g44169 not n15644 ; n15644_not
g44170 not n15635 ; n15635_not
g44171 not n17642 ; n17642_not
g44172 not n15626 ; n15626_not
g44173 not n17651 ; n17651_not
g44174 not n15617 ; n15617_not
g44175 not n18551 ; n18551_not
g44176 not n11963 ; n11963_not
g44177 not n25562 ; n25562_not
g44178 not n25508 ; n25508_not
g44179 not n25634 ; n25634_not
g44180 not n25643 ; n25643_not
g44181 not n11954 ; n11954_not
g44182 not n25652 ; n25652_not
g44183 not n19280 ; n19280_not
g44184 not n25661 ; n25661_not
g44185 not n25670 ; n25670_not
g44186 not n11891 ; n11891_not
g44187 not n11945 ; n11945_not
g44188 not n25706 ; n25706_not
g44189 not n19262 ; n19262_not
g44190 not n11936 ; n11936_not
g44191 not n25625 ; n25625_not
g44192 not n11927 ; n11927_not
g44193 not n19253 ; n19253_not
g44194 not n25733 ; n25733_not
g44195 not n18380 ; n18380_not
g44196 not n11909 ; n11909_not
g44197 not n25517 ; n25517_not
g44198 not n12098 ; n12098_not
g44199 not n12089 ; n12089_not
g44200 not n19334 ; n19334_not
g44201 not n25526 ; n25526_not
g44202 not n18416 ; n18416_not
g44203 not n19325 ; n19325_not
g44204 not n11855 ; n11855_not
g44205 not n11657 ; n11657_not
g44206 not n18542 ; n18542_not
g44207 not n19316 ; n19316_not
g44208 not n25544 ; n25544_not
g44209 not n25553 ; n25553_not
g44210 not n11990 ; n11990_not
g44211 not n25463 ; n25463_not
g44212 not n19307 ; n19307_not
g44213 not n11981 ; n11981_not
g44214 not n25571 ; n25571_not
g44215 not n25580 ; n25580_not
g44216 not n25607 ; n25607_not
g44217 not n19019 ; n19019_not
g44218 not n11972 ; n11972_not
g44219 not n25616 ; n25616_not
g44220 not n19190 ; n19190_not
g44221 not n11783 ; n11783_not
g44222 not n11837 ; n11837_not
g44223 not n11819 ; n11819_not
g44224 not n19172 ; n19172_not
g44225 not n11792 ; n11792_not
g44226 not n26039 ; n26039_not
g44227 not n26057 ; n26057_not
g44228 not n19163 ; n19163_not
g44229 not n19154 ; n19154_not
g44230 not n11747 ; n11747_not
g44231 not n26075 ; n26075_not
g44232 not n11738 ; n11738_not
g44233 not n11729 ; n11729_not
g44234 not n26084 ; n26084_not
g44235 not n19145 ; n19145_not
g44236 not n26066 ; n26066_not
g44237 not n26093 ; n26093_not
g44238 not n11684 ; n11684_not
g44239 not n11675 ; n11675_not
g44240 not n11666 ; n11666_not
g44241 not n19127 ; n19127_not
g44242 not n11648 ; n11648_not
g44243 not n19118 ; n19118_not
g44244 not n19244 ; n19244_not
g44245 not n11918 ; n11918_not
g44246 not n25742 ; n25742_not
g44247 not n25751 ; n25751_not
g44248 not n19235 ; n19235_not
g44249 not n18560 ; n18560_not
g44250 not n25760 ; n25760_not
g44251 not n19226 ; n19226_not
g44252 not n25814 ; n25814_not
g44253 not n11882 ; n11882_not
g44254 not n25823 ; n25823_not
g44255 not n25805 ; n25805_not
g44256 not n19217 ; n19217_not
g44257 not n25841 ; n25841_not
g44258 not n25850 ; n25850_not
g44259 not n19208 ; n19208_not
g44260 not n11864 ; n11864_not
g44261 not n25913 ; n25913_not
g44262 not n25922 ; n25922_not
g44263 not n25931 ; n25931_not
g44264 not n11594 ; n11594_not
g44265 not n25940 ; n25940_not
g44266 not n19514 ; n19514_not
g44267 not n12674 ; n12674_not
g44268 not n19523 ; n19523_not
g44269 not n25238 ; n25238_not
g44270 not n12665 ; n12665_not
g44271 not n25247 ; n25247_not
g44272 not n19136 ; n19136_not
g44273 not n12656 ; n12656_not
g44274 not n25256 ; n25256_not
g44275 not n19505 ; n19505_not
g44276 not n25076 ; n25076_not
g44277 not n12629 ; n12629_not
g44278 not n25265 ; n25265_not
g44279 not n25274 ; n25274_not
g44280 not n25283 ; n25283_not
g44281 not n12593 ; n12593_not
g44282 not n12197 ; n12197_not
g44283 not n12575 ; n12575_not
g44284 not n12566 ; n12566_not
g44285 not n25319 ; n25319_not
g44286 not n19460 ; n19460_not
g44287 not n12557 ; n12557_not
g44288 not n12548 ; n12548_not
g44289 not n12539 ; n12539_not
g44290 not n12827 ; n12827_not
g44291 not n12809 ; n12809_not
g44292 not n24950 ; n24950_not
g44293 not n18470 ; n18470_not
g44294 not n12791 ; n12791_not
g44295 not n25139 ; n25139_not
g44296 not n12782 ; n12782_not
g44297 not n24626 ; n24626_not
g44298 not n25148 ; n25148_not
g44299 not n12773 ; n12773_not
g44300 not n25157 ; n25157_not
g44301 not n12764 ; n12764_not
g44302 not n25166 ; n25166_not
g44303 not n25175 ; n25175_not
g44304 not n25184 ; n25184_not
g44305 not n19550 ; n19550_not
g44306 not n12746 ; n12746_not
g44307 not n25193 ; n25193_not
g44308 not n19541 ; n19541_not
g44309 not n12737 ; n12737_not
g44310 not n12719 ; n12719_not
g44311 not n12728 ; n12728_not
g44312 not n12683 ; n12683_not
g44313 not n12647 ; n12647_not
g44314 not n25229 ; n25229_not
g44315 not n25409 ; n25409_not
g44316 not n25328 ; n25328_not
g44317 not n12386 ; n12386_not
g44318 not n12377 ; n12377_not
g44319 not n12368 ; n12368_not
g44320 not n12359 ; n12359_not
g44321 not n25427 ; n25427_not
g44322 not n25436 ; n25436_not
g44323 not n25445 ; n25445_not
g44324 not n25292 ; n25292_not
g44325 not n19370 ; n19370_not
g44326 not n25454 ; n25454_not
g44327 not n12287 ; n12287_not
g44328 not n12269 ; n12269_not
g44329 not n25472 ; n25472_not
g44330 not n25490 ; n25490_not
g44331 not n19343 ; n19343_not
g44332 not n19352 ; n19352_not
g44333 not n12188 ; n12188_not
g44334 not n18533 ; n18533_not
g44335 not n11828 ; n11828_not
g44336 not n25337 ; n25337_not
g44337 not n12278 ; n12278_not
g44338 not n25346 ; n25346_not
g44339 not n19451 ; n19451_not
g44340 not n12494 ; n12494_not
g44341 not n12485 ; n12485_not
g44342 not n19442 ; n19442_not
g44343 not n25355 ; n25355_not
g44344 not n12476 ; n12476_not
g44345 not n25364 ; n25364_not
g44346 not n12467 ; n12467_not
g44347 not n25382 ; n25382_not
g44348 not n25391 ; n25391_not
g44349 not n19424 ; n19424_not
g44350 not n18506 ; n18506_not
g44351 not n12458 ; n12458_not
g44352 not n19415 ; n19415_not
g44353 not n12449 ; n12449_not
g44354 not n18515 ; n18515_not
g44355 not n19406 ; n19406_not
g44356 not n18524 ; n18524_not
g44357 not n12395 ; n12395_not
g44358 not n26660 ; n26660_not
g44359 not n10685 ; n10685_not
g44360 not n26633 ; n26633_not
g44361 not n26705 ; n26705_not
g44362 not n10667 ; n10667_not
g44363 not n10658 ; n10658_not
g44364 not n10649 ; n10649_not
g44365 not n26723 ; n26723_not
g44366 not n26714 ; n26714_not
g44367 not n26732 ; n26732_not
g44368 not n26741 ; n26741_not
g44369 not n26750 ; n26750_not
g44370 not n18830 ; n18830_not
g44371 not n26804 ; n26804_not
g44372 not n10595 ; n10595_not
g44373 not n10586 ; n10586_not
g44374 not n26813 ; n26813_not
g44375 not n18821 ; n18821_not
g44376 not n10577 ; n10577_not
g44377 not n26822 ; n26822_not
g44378 not n26831 ; n26831_not
g44379 not n18812 ; n18812_not
g44380 not n10568 ; n10568_not
g44381 not n10559 ; n10559_not
g44382 not n26903 ; n26903_not
g44383 not n26507 ; n26507_not
g44384 not n10793 ; n10793_not
g44385 not n18911 ; n18911_not
g44386 not n26525 ; n26525_not
g44387 not n26516 ; n26516_not
g44388 not n10775 ; n10775_not
g44389 not n26534 ; n26534_not
g44390 not n26453 ; n26453_not
g44391 not n26543 ; n26543_not
g44392 not n10766 ; n10766_not
g44393 not n26552 ; n26552_not
g44394 not n10757 ; n10757_not
g44395 not n26561 ; n26561_not
g44396 not n26570 ; n26570_not
g44397 not n10469 ; n10469_not
g44398 not n10748 ; n10748_not
g44399 not n26606 ; n26606_not
g44400 not n10739 ; n10739_not
g44401 not n10694 ; n10694_not
g44402 not n26615 ; n26615_not
g44403 not n26642 ; n26642_not
g44404 not n18722 ; n18722_not
g44405 not n18731 ; n18731_not
g44406 not n27146 ; n27146_not
g44407 not n27128 ; n27128_not
g44408 not n27155 ; n27155_not
g44409 not n27164 ; n27164_not
g44410 not n27173 ; n27173_not
g44411 not n27182 ; n27182_not
g44412 not n27191 ; n27191_not
g44413 not n27209 ; n27209_not
g44414 not n18713 ; n18713_not
g44415 not n27218 ; n27218_not
g44416 not n27227 ; n27227_not
g44417 not n27245 ; n27245_not
g44418 not n18704 ; n18704_not
g44419 not n27254 ; n27254_not
g44420 not n27263 ; n27263_not
g44421 not n27272 ; n27272_not
g44422 not n27281 ; n27281_not
g44423 not n27308 ; n27308_not
g44424 not n27317 ; n27317_not
g44425 not n26840 ; n26840_not
g44426 not n26912 ; n26912_not
g44427 not n10199 ; n10199_not
g44428 not n26921 ; n26921_not
g44429 not n26930 ; n26930_not
g44430 not n10496 ; n10496_not
g44431 not n10478 ; n10478_not
g44432 not n10379 ; n10379_not
g44433 not n10388 ; n10388_not
g44434 not n10298 ; n10298_not
g44435 not n27029 ; n27029_not
g44436 not n10289 ; n10289_not
g44437 not n27038 ; n27038_not
g44438 not n27056 ; n27056_not
g44439 not n27065 ; n27065_not
g44440 not n27074 ; n27074_not
g44441 not n27119 ; n27119_not
g44442 not n27137 ; n27137_not
g44443 not n19073 ; n19073_not
g44444 not n11387 ; n11387_not
g44445 not n11396 ; n11396_not
g44446 not n11378 ; n11378_not
g44447 not n18335 ; n18335_not
g44448 not n11369 ; n11369_not
g44449 not n26219 ; n26219_not
g44450 not n19055 ; n19055_not
g44451 not n18632 ; n18632_not
g44452 not n11297 ; n11297_not
g44453 not n19046 ; n19046_not
g44454 not n11288 ; n11288_not
g44455 not n26228 ; n26228_not
g44456 not n11279 ; n11279_not
g44457 not n18641 ; n18641_not
g44458 not n11189 ; n11189_not
g44459 not n19037 ; n19037_not
g44460 not n11198 ; n11198_not
g44461 not n26237 ; n26237_not
g44462 not n19028 ; n19028_not
g44463 not n10847 ; n10847_not
g44464 not n10856 ; n10856_not
g44465 not n18605 ; n18605_not
g44466 not n26129 ; n26129_not
g44467 not n11585 ; n11585_not
g44468 not n19109 ; n19109_not
g44469 not n18614 ; n18614_not
g44470 not n11576 ; n11576_not
g44471 not n18623 ; n18623_not
g44472 not n26138 ; n26138_not
g44473 not n11558 ; n11558_not
g44474 not n26147 ; n26147_not
g44475 not n11495 ; n11495_not
g44476 not n19091 ; n19091_not
g44477 not n11549 ; n11549_not
g44478 not n26165 ; n26165_not
g44479 not n19082 ; n19082_not
g44480 not n26174 ; n26174_not
g44481 not n11486 ; n11486_not
g44482 not n26183 ; n26183_not
g44483 not n11477 ; n11477_not
g44484 not n11468 ; n11468_not
g44485 not n10919 ; n10919_not
g44486 not n26363 ; n26363_not
g44487 not n26372 ; n26372_not
g44488 not n26381 ; n26381_not
g44489 not n26390 ; n26390_not
g44490 not n10892 ; n10892_not
g44491 not n10883 ; n10883_not
g44492 not n26408 ; n26408_not
g44493 not n10487 ; n10487_not
g44494 not n26417 ; n26417_not
g44495 not n26318 ; n26318_not
g44496 not n10874 ; n10874_not
g44497 not n26426 ; n26426_not
g44498 not n10865 ; n10865_not
g44499 not n26435 ; n26435_not
g44500 not n26444 ; n26444_not
g44501 not n26462 ; n26462_not
g44502 not n26471 ; n26471_not
g44503 not n26480 ; n26480_not
g44504 not n10838 ; n10838_not
g44505 not n10829 ; n10829_not
g44506 not n18650 ; n18650_not
g44507 not n26246 ; n26246_not
g44508 not n10982 ; n10982_not
g44509 not n26255 ; n26255_not
g44510 not n26264 ; n26264_not
g44511 not n18317 ; n18317_not
g44512 not n26273 ; n26273_not
g44513 not n10991 ; n10991_not
g44514 not n26282 ; n26282_not
g44515 not n26309 ; n26309_not
g44516 not n10973 ; n10973_not
g44517 not n10964 ; n10964_not
g44518 not n26327 ; n26327_not
g44519 not n26336 ; n26336_not
g44520 not n10946 ; n10946_not
g44521 not n10937 ; n10937_not
g44522 not n26345 ; n26345_not
g44523 not n10928 ; n10928_not
g44524 not n26354 ; n26354_not
g44525 not n19901 ; n19901_not
g44526 not n24671 ; n24671_not
g44527 not n24932 ; n24932_not
g44528 not n13538 ; n13538_not
g44529 not n19721 ; n19721_not
g44530 not n19820 ; n19820_not
g44531 not n13754 ; n13754_not
g44532 not n24491 ; n24491_not
g44533 not n24923 ; n24923_not
g44534 not n24329 ; n24329_not
g44535 not n19631 ; n19631_not
g44536 not n24680 ; n24680_not
g44537 not n13736 ; n13736_not
g44538 not n24914 ; n24914_not
g44539 not n18443 ; n18443_not
g44540 not n12980 ; n12980_not
g44541 not n13727 ; n13727_not
g44542 not n19640 ; n19640_not
g44543 not n13196 ; n13196_not
g44544 not n13718 ; n13718_not
g44545 not n24473 ; n24473_not
g44546 not n12944 ; n12944_not
g44547 not n24275 ; n24275_not
g44548 not n13781 ; n13781_not
g44549 not n12953 ; n12953_not
g44550 not n13259 ; n13259_not
g44551 not n19622 ; n19622_not
g44552 not n18461 ; n18461_not
g44553 not n24284 ; n24284_not
g44554 not n24518 ; n24518_not
g44555 not n12971 ; n12971_not
g44556 not n24653 ; n24653_not
g44557 not n24293 ; n24293_not
g44558 not n24464 ; n24464_not
g44559 not n24509 ; n24509_not
g44560 not n19730 ; n19730_not
g44561 not n13493 ; n13493_not
g44562 not n24662 ; n24662_not
g44563 not n13772 ; n13772_not
g44564 not n19613 ; n19613_not
g44565 not n24941 ; n24941_not
g44566 not n24257 ; n24257_not
g44567 not n24383 ; n24383_not
g44568 not n13574 ; n13574_not
g44569 not n24770 ; n24770_not
g44570 not n24590 ; n24590_not
g44571 not n13646 ; n13646_not
g44572 not n24455 ; n24455_not
g44573 not n12755 ; n12755_not
g44574 not n24761 ; n24761_not
g44575 not n24725 ; n24725_not
g44576 not n24752 ; n24752_not
g44577 not n13628 ; n13628_not
g44578 not n13619 ; n13619_not
g44579 not n24428 ; n24428_not
g44580 not n24743 ; n24743_not
g44581 not n13097 ; n13097_not
g44582 not n13079 ; n13079_not
g44583 not n24437 ; n24437_not
g44584 not n13583 ; n13583_not
g44585 not n24734 ; n24734_not
g44586 not n24446 ; n24446_not
g44587 not n13088 ; n13088_not
g44588 not n13187 ; n13187_not
g44589 not n24707 ; n24707_not
g44590 not n13709 ; n13709_not
g44591 not n24860 ; n24860_not
g44592 not n24347 ; n24347_not
g44593 not n24851 ; n24851_not
g44594 not n19712 ; n19712_not
g44595 not n24338 ; n24338_not
g44596 not n24833 ; n24833_not
g44597 not n24842 ; n24842_not
g44598 not n13178 ; n13178_not
g44599 not n24482 ; n24482_not
g44600 not n13565 ; n13565_not
g44601 not n24824 ; n24824_not
g44602 not n19703 ; n19703_not
g44603 not n24356 ; n24356_not
g44604 not n13682 ; n13682_not
g44605 not n13169 ; n13169_not
g44606 not n24365 ; n24365_not
g44607 not n24815 ; n24815_not
g44608 not n18452 ; n18452_not
g44609 not n24716 ; n24716_not
g44610 not n24806 ; n24806_not
g44611 not n25067 ; n25067_not
g44612 not n13277 ; n13277_not
g44613 not n24266 ; n24266_not
g44614 not n24545 ; n24545_not
g44615 not n13835 ; n13835_not
g44616 not n25049 ; n25049_not
g44617 not n13448 ; n13448_not
g44618 not n13457 ; n13457_not
g44619 not n13394 ; n13394_not
g44620 not n13358 ; n13358_not
g44621 not n25094 ; n25094_not
g44622 not n13286 ; n13286_not
g44623 not n12863 ; n12863_not
g44624 not n24635 ; n24635_not
g44625 not n24239 ; n24239_not
g44626 not n13439 ; n13439_not
g44627 not n13817 ; n13817_not
g44628 not n13871 ; n13871_not
g44629 not n24563 ; n24563_not
g44630 not n13367 ; n13367_not
g44631 not n25058 ; n25058_not
g44632 not n13349 ; n13349_not
g44633 not n12890 ; n12890_not
g44634 not n19604 ; n19604_not
g44635 not n24608 ; n24608_not
g44636 not n12881 ; n12881_not
g44637 not n13880 ; n13880_not
g44638 not n12845 ; n12845_not
g44639 not n13853 ; n13853_not
g44640 not n24554 ; n24554_not
g44641 not n13475 ; n13475_not
g44642 not n24527 ; n24527_not
g44643 not n13268 ; n13268_not
g44644 not n19802 ; n19802_not
g44645 not n12926 ; n12926_not
g44646 not n12917 ; n12917_not
g44647 not n25085 ; n25085_not
g44648 not n13376 ; n13376_not
g44649 not n12908 ; n12908_not
g44650 not n13295 ; n13295_not
g44651 not n24581 ; n24581_not
g44652 not n24194 ; n24194_not
g44653 not n24536 ; n24536_not
g44654 not n13484 ; n13484_not
g44655 not n23907 ; n23907_not
g44656 not n16455 ; n16455_not
g44657 not n23754 ; n23754_not
g44658 not n21963 ; n21963_not
g44659 not n16095 ; n16095_not
g44660 not n21954 ; n21954_not
g44661 not n10884 ; n10884_not
g44662 not n13566 ; n13566_not
g44663 not n26166 ; n26166_not
g44664 not n10866 ; n10866_not
g44665 not n16077 ; n16077_not
g44666 not n26391 ; n26391_not
g44667 not n24465 ; n24465_not
g44668 not n10893 ; n10893_not
g44669 not n14457 ; n14457_not
g44670 not n16086 ; n16086_not
g44671 not n11496 ; n11496_not
g44672 not n21729 ; n21729_not
g44673 not n11487 ; n11487_not
g44674 not n22188 ; n22188_not
g44675 not n13557 ; n13557_not
g44676 not n23709 ; n23709_not
g44677 not n13395 ; n13395_not
g44678 not n21972 ; n21972_not
g44679 not n26409 ; n26409_not
g44680 not n13296 ; n13296_not
g44681 not n14448 ; n14448_not
g44682 not n21990 ; n21990_not
g44683 not n26355 ; n26355_not
g44684 not n21918 ; n21918_not
g44685 not n24438 ; n24438_not
g44686 not n26418 ; n26418_not
g44687 not n16059 ; n16059_not
g44688 not n26445 ; n26445_not
g44689 not n26148 ; n26148_not
g44690 not n24447 ; n24447_not
g44691 not n10767 ; n10767_not
g44692 not n24573 ; n24573_not
g44693 not n14475 ; n14475_not
g44694 not n10857 ; n10857_not
g44695 not n11559 ; n11559_not
g44696 not n15627 ; n15627_not
g44697 not n26139 ; n26139_not
g44698 not n23925 ; n23925_not
g44699 not n23745 ; n23745_not
g44700 not n14286 ; n14286_not
g44701 not n16482 ; n16482_not
g44702 not n21909 ; n21909_not
g44703 not n26454 ; n26454_not
g44704 not n15960 ; n15960_not
g44705 not n26463 ; n26463_not
g44706 not n16446 ; n16446_not
g44707 not n13575 ; n13575_not
g44708 not n10875 ; n10875_not
g44709 not n23916 ; n23916_not
g44710 not n24564 ; n24564_not
g44711 not n21945 ; n21945_not
g44712 not n16464 ; n16464_not
g44713 not n21936 ; n21936_not
g44714 not n14295 ; n14295_not
g44715 not n16068 ; n16068_not
g44716 not n13449 ; n13449_not
g44717 not n14277 ; n14277_not
g44718 not n26436 ; n26436_not
g44719 not n16473 ; n16473_not
g44720 not n21927 ; n21927_not
g44721 not n14466 ; n14466_not
g44722 not n16266 ; n16266_not
g44723 not n26427 ; n26427_not
g44724 not n16167 ; n16167_not
g44725 not n26256 ; n26256_not
g44726 not n13458 ; n13458_not
g44727 not n11298 ; n11298_not
g44728 not n26265 ; n26265_not
g44729 not n13485 ; n13485_not
g44730 not n23835 ; n23835_not
g44731 not n10992 ; n10992_not
g44732 not n16275 ; n16275_not
g44733 not n23682 ; n23682_not
g44734 not n26283 ; n26283_not
g44735 not n16284 ; n16284_not
g44736 not n16293 ; n16293_not
g44737 not n23790 ; n23790_not
g44738 not n22089 ; n22089_not
g44739 not n10983 ; n10983_not
g44740 not n24546 ; n24546_not
g44741 not n13539 ; n13539_not
g44742 not n16329 ; n16329_not
g44743 not n23781 ; n23781_not
g44744 not n26238 ; n26238_not
g44745 not n15861 ; n15861_not
g44746 not n14394 ; n14394_not
g44747 not n23808 ; n23808_not
g44748 not n16239 ; n16239_not
g44749 not n24519 ; n24519_not
g44750 not n11199 ; n11199_not
g44751 not n14385 ; n14385_not
g44752 not n16194 ; n16194_not
g44753 not n13476 ; n13476_not
g44754 not n16185 ; n16185_not
g44755 not n16248 ; n16248_not
g44756 not n26247 ; n26247_not
g44757 not n13098 ; n13098_not
g44758 not n23826 ; n23826_not
g44759 not n24528 ; n24528_not
g44760 not n16257 ; n16257_not
g44761 not n13467 ; n13467_not
g44762 not n13494 ; n13494_not
g44763 not n16176 ; n16176_not
g44764 not n14439 ; n14439_not
g44765 not n11289 ; n11289_not
g44766 not n24537 ; n24537_not
g44767 not n10938 ; n10938_not
g44768 not n15816 ; n15816_not
g44769 not n15951 ; n15951_not
g44770 not n11469 ; n11469_not
g44771 not n23880 ; n23880_not
g44772 not n26346 ; n26346_not
g44773 not n26193 ; n26193_not
g44774 not n10929 ; n10929_not
g44775 not n22179 ; n22179_not
g44776 not n24483 ; n24483_not
g44777 not n14349 ; n14349_not
g44778 not n23772 ; n23772_not
g44779 not n24555 ; n24555_not
g44780 not n26184 ; n26184_not
g44781 not n26274 ; n26274_not
g44782 not n16419 ; n16419_not
g44783 not n16428 ; n16428_not
g44784 not n23763 ; n23763_not
g44785 not n24474 ; n24474_not
g44786 not n26364 ; n26364_not
g44787 not n16437 ; n16437_not
g44788 not n14367 ; n14367_not
g44789 not n11379 ; n11379_not
g44790 not n16338 ; n16338_not
g44791 not n26319 ; n26319_not
g44792 not n10965 ; n10965_not
g44793 not n23853 ; n23853_not
g44794 not n11397 ; n11397_not
g44795 not n16347 ; n16347_not
g44796 not n16356 ; n16356_not
g44797 not n10947 ; n10947_not
g44798 not n21981 ; n21981_not
g44799 not n13548 ; n13548_not
g44800 not n16365 ; n16365_not
g44801 not n26175 ; n26175_not
g44802 not n26337 ; n26337_not
g44803 not n26328 ; n26328_not
g44804 not n13278 ; n13278_not
g44805 not n23862 ; n23862_not
g44806 not n16383 ; n16383_not
g44807 not n13782 ; n13782_not
g44808 not n10299 ; n10299_not
g44809 not n24087 ; n24087_not
g44810 not n21567 ; n21567_not
g44811 not n24096 ; n24096_not
g44812 not n13980 ; n13980_not
g44813 not n16770 ; n16770_not
g44814 not n21558 ; n21558_not
g44815 not n27039 ; n27039_not
g44816 not n13971 ; n13971_not
g44817 not n27057 ; n27057_not
g44818 not n21549 ; n21549_not
g44819 not n27048 ; n27048_not
g44820 not n13890 ; n13890_not
g44821 not n27066 ; n27066_not
g44822 not n24267 ; n24267_not
g44823 not n27075 ; n27075_not
g44824 not n27084 ; n27084_not
g44825 not n27093 ; n27093_not
g44826 not n16806 ; n16806_not
g44827 not n27129 ; n27129_not
g44828 not n13962 ; n13962_not
g44829 not n26832 ; n26832_not
g44830 not n13845 ; n13845_not
g44831 not n26850 ; n26850_not
g44832 not n14097 ; n14097_not
g44833 not n13368 ; n13368_not
g44834 not n21459 ; n21459_not
g44835 not n26904 ; n26904_not
g44836 not n26841 ; n26841_not
g44837 not n13773 ; n13773_not
g44838 not n16725 ; n16725_not
g44839 not n14088 ; n14088_not
g44840 not n26913 ; n26913_not
g44841 not n16734 ; n16734_not
g44842 not n10389 ; n10389_not
g44843 not n21585 ; n21585_not
g44844 not n10398 ; n10398_not
g44845 not n16743 ; n16743_not
g44846 not n14079 ; n14079_not
g44847 not n10479 ; n10479_not
g44848 not n16752 ; n16752_not
g44849 not n10488 ; n10488_not
g44850 not n10497 ; n10497_not
g44851 not n24069 ; n24069_not
g44852 not n26940 ; n26940_not
g44853 not n26931 ; n26931_not
g44854 not n26922 ; n26922_not
g44855 not n24294 ; n24294_not
g44856 not n13917 ; n13917_not
g44857 not n16860 ; n16860_not
g44858 not n16518 ; n16518_not
g44859 not n13863 ; n13863_not
g44860 not n16905 ; n16905_not
g44861 not n21396 ; n21396_not
g44862 not n13881 ; n13881_not
g44863 not n27255 ; n27255_not
g44864 not n27246 ; n27246_not
g44865 not n27237 ; n27237_not
g44866 not n24195 ; n24195_not
g44867 not n16923 ; n16923_not
g44868 not n21378 ; n21378_not
g44869 not n13908 ; n13908_not
g44870 not n27273 ; n27273_not
g44871 not n16932 ; n16932_not
g44872 not n27282 ; n27282_not
g44873 not n16545 ; n16545_not
g44874 not n21369 ; n21369_not
g44875 not n16833 ; n16833_not
g44876 not n16941 ; n16941_not
g44877 not n27291 ; n27291_not
g44878 not n24177 ; n24177_not
g44879 not n16950 ; n16950_not
g44880 not n24186 ; n24186_not
g44881 not n27138 ; n27138_not
g44882 not n24258 ; n24258_not
g44883 not n13719 ; n13719_not
g44884 not n27147 ; n27147_not
g44885 not n13953 ; n13953_not
g44886 not n16824 ; n16824_not
g44887 not n21486 ; n21486_not
g44888 not n27156 ; n27156_not
g44889 not n13818 ; n13818_not
g44890 not n13944 ; n13944_not
g44891 not n21495 ; n21495_not
g44892 not n27174 ; n27174_not
g44893 not n13827 ; n13827_not
g44894 not n27183 ; n27183_not
g44895 not n27219 ; n27219_not
g44896 not n24159 ; n24159_not
g44897 not n16851 ; n16851_not
g44898 not n21468 ; n21468_not
g44899 not n13854 ; n13854_not
g44900 not n13926 ; n13926_not
g44901 not n27165 ; n27165_not
g44902 not n27192 ; n27192_not
g44903 not n16842 ; n16842_not
g44904 not n13836 ; n13836_not
g44905 not n13935 ; n13935_not
g44906 not n13638 ; n13638_not
g44907 not n26553 ; n26553_not
g44908 not n14259 ; n14259_not
g44909 not n13656 ; n13656_not
g44910 not n26562 ; n26562_not
g44911 not n24384 ; n24384_not
g44912 not n16554 ; n16554_not
g44913 not n26571 ; n26571_not
g44914 not n10758 ; n10758_not
g44915 not n16563 ; n16563_not
g44916 not n10749 ; n10749_not
g44917 not n13674 ; n13674_not
g44918 not n24375 ; n24375_not
g44919 not n16572 ; n16572_not
g44920 not n21792 ; n21792_not
g44921 not n24366 ; n24366_not
g44922 not n26616 ; n26616_not
g44923 not n10695 ; n10695_not
g44924 not n21783 ; n21783_not
g44925 not n24357 ; n24357_not
g44926 not n16581 ; n16581_not
g44927 not n26625 ; n26625_not
g44928 not n21765 ; n21765_not
g44929 not n26382 ; n26382_not
g44930 not n16491 ; n16491_not
g44931 not n26472 ; n26472_not
g44932 not n26481 ; n26481_not
g44933 not n10848 ; n10848_not
g44934 not n21864 ; n21864_not
g44935 not n10839 ; n10839_not
g44936 not n16509 ; n16509_not
g44937 not n24429 ; n24429_not
g44938 not n21855 ; n21855_not
g44939 not n13593 ; n13593_not
g44940 not n26508 ; n26508_not
g44941 not n26544 ; n26544_not
g44942 not n14268 ; n14268_not
g44943 not n21828 ; n21828_not
g44944 not n10776 ; n10776_not
g44945 not n26535 ; n26535_not
g44946 not n23970 ; n23970_not
g44947 not n16527 ; n16527_not
g44948 not n21846 ; n21846_not
g44949 not n13629 ; n13629_not
g44950 not n26490 ; n26490_not
g44951 not n23961 ; n23961_not
g44952 not n26526 ; n26526_not
g44953 not n26517 ; n26517_not
g44954 not n10794 ; n10794_not
g44955 not n26733 ; n26733_not
g44956 not n13728 ; n13728_not
g44957 not n16653 ; n16653_not
g44958 not n26742 ; n26742_not
g44959 not n16662 ; n16662_not
g44960 not n21693 ; n21693_not
g44961 not n14169 ; n14169_not
g44962 not n26751 ; n26751_not
g44963 not n26760 ; n26760_not
g44964 not n10596 ; n10596_not
g44965 not n13737 ; n13737_not
g44966 not n21684 ; n21684_not
g44967 not n13755 ; n13755_not
g44968 not n26823 ; n26823_not
g44969 not n16707 ; n16707_not
g44970 not n13809 ; n13809_not
g44971 not n21639 ; n21639_not
g44972 not n10578 ; n10578_not
g44973 not n21648 ; n21648_not
g44974 not n21387 ; n21387_not
g44975 not n26814 ; n26814_not
g44976 not n16680 ; n16680_not
g44977 not n16671 ; n16671_not
g44978 not n10587 ; n10587_not
g44979 not n21675 ; n21675_not
g44980 not n16590 ; n16590_not
g44981 not n14196 ; n14196_not
g44982 not n21747 ; n21747_not
g44983 not n13692 ; n13692_not
g44984 not n26634 ; n26634_not
g44985 not n10686 ; n10686_not
g44986 not n13791 ; n13791_not
g44987 not n16617 ; n16617_not
g44988 not n26580 ; n26580_not
g44989 not n26643 ; n26643_not
g44990 not n26652 ; n26652_not
g44991 not n14187 ; n14187_not
g44992 not n26661 ; n26661_not
g44993 not n26706 ; n26706_not
g44994 not n26724 ; n26724_not
g44995 not n16644 ; n16644_not
g44996 not n14178 ; n14178_not
g44997 not n26715 ; n26715_not
g44998 not n24339 ; n24339_not
g44999 not n10659 ; n10659_not
g45000 not n16635 ; n16635_not
g45001 not n10668 ; n10668_not
g45002 not n24348 ; n24348_not
g45003 not n16626 ; n16626_not
g45004 not n26670 ; n26670_not
g45005 not n25392 ; n25392_not
g45006 not n15276 ; n15276_not
g45007 not n24924 ; n24924_not
g45008 not n15285 ; n15285_not
g45009 not n24915 ; n24915_not
g45010 not n15294 ; n15294_not
g45011 not n22782 ; n22782_not
g45012 not n14655 ; n14655_not
g45013 not n12396 ; n12396_not
g45014 not n25329 ; n25329_not
g45015 not n23538 ; n23538_not
g45016 not n15339 ; n15339_not
g45017 not n23547 ; n23547_not
g45018 not n25428 ; n25428_not
g45019 not n22971 ; n22971_not
g45020 not n24906 ; n24906_not
g45021 not n25257 ; n25257_not
g45022 not n12369 ; n12369_not
g45023 not n25419 ; n25419_not
g45024 not n15375 ; n15375_not
g45025 not n12378 ; n12378_not
g45026 not n15357 ; n15357_not
g45027 not n12981 ; n12981_not
g45028 not n12387 ; n12387_not
g45029 not n14961 ; n14961_not
g45030 not n15348 ; n15348_not
g45031 not n14646 ; n14646_not
g45032 not n15177 ; n15177_not
g45033 not n23097 ; n23097_not
g45034 not n25347 ; n25347_not
g45035 not n12495 ; n12495_not
g45036 not n24942 ; n24942_not
g45037 not n23088 ; n23088_not
g45038 not n14673 ; n14673_not
g45039 not n15195 ; n15195_not
g45040 not n12486 ; n12486_not
g45041 not n22818 ; n22818_not
g45042 not n12279 ; n12279_not
g45043 not n25356 ; n25356_not
g45044 not n23079 ; n23079_not
g45045 not n22980 ; n22980_not
g45046 not n23529 ; n23529_not
g45047 not n24735 ; n24735_not
g45048 not n25383 ; n25383_not
g45049 not n12459 ; n12459_not
g45050 not n15267 ; n15267_not
g45051 not n14664 ; n14664_not
g45052 not n15258 ; n15258_not
g45053 not n25374 ; n25374_not
g45054 not n12468 ; n12468_not
g45055 not n24933 ; n24933_not
g45056 not n25365 ; n25365_not
g45057 not n15249 ; n15249_not
g45058 not n12189 ; n12189_not
g45059 not n24690 ; n24690_not
g45060 not n22890 ; n22890_not
g45061 not n15447 ; n15447_not
g45062 not n22881 ; n22881_not
g45063 not n24816 ; n24816_not
g45064 not n22872 ; n22872_not
g45065 not n22863 ; n22863_not
g45066 not n22854 ; n22854_not
g45067 not n15456 ; n15456_not
g45068 not n25509 ; n25509_not
g45069 not n23565 ; n23565_not
g45070 not n22845 ; n22845_not
g45071 not n25527 ; n25527_not
g45072 not n15483 ; n15483_not
g45073 not n23583 ; n23583_not
g45074 not n24780 ; n24780_not
g45075 not n22827 ; n22827_not
g45076 not n12684 ; n12684_not
g45077 not n12693 ; n12693_not
g45078 not n12099 ; n12099_not
g45079 not n25518 ; n25518_not
g45080 not n22836 ; n22836_not
g45081 not n15465 ; n15465_not
g45082 not n24807 ; n24807_not
g45083 not n15393 ; n15393_not
g45084 not n24843 ; n24843_not
g45085 not n23556 ; n23556_not
g45086 not n22935 ; n22935_not
g45087 not n22944 ; n22944_not
g45088 not n15384 ; n15384_not
g45089 not n25446 ; n25446_not
g45090 not n25293 ; n25293_not
g45091 not n22953 ; n22953_not
g45092 not n22962 ; n22962_not
g45093 not n25437 ; n25437_not
g45094 not n24861 ; n24861_not
g45095 not n12927 ; n12927_not
g45096 not n15438 ; n15438_not
g45097 not n15429 ; n15429_not
g45098 not n24825 ; n24825_not
g45099 not n12198 ; n12198_not
g45100 not n23574 ; n23574_not
g45101 not n25491 ; n25491_not
g45102 not n25482 ; n25482_not
g45103 not n25473 ; n25473_not
g45104 not n14619 ; n14619_not
g45105 not n22908 ; n22908_not
g45106 not n24834 ; n24834_not
g45107 not n25464 ; n25464_not
g45108 not n14628 ; n14628_not
g45109 not n12288 ; n12288_not
g45110 not n22917 ; n22917_not
g45111 not n25095 ; n25095_not
g45112 not n25167 ; n25167_not
g45113 not n25176 ; n25176_not
g45114 not n25086 ; n25086_not
g45115 not n14853 ; n14853_not
g45116 not n12756 ; n12756_not
g45117 not n12738 ; n12738_not
g45118 not n12747 ; n12747_not
g45119 not n14862 ; n14862_not
g45120 not n14763 ; n14763_not
g45121 not n14871 ; n14871_not
g45122 not n25185 ; n25185_not
g45123 not n14880 ; n14880_not
g45124 not n12864 ; n12864_not
g45125 not n12882 ; n12882_not
g45126 not n23268 ; n23268_not
g45127 not n14745 ; n14745_not
g45128 not n14907 ; n14907_not
g45129 not n23448 ; n23448_not
g45130 not n12729 ; n12729_not
g45131 not n23439 ; n23439_not
g45132 not n23277 ; n23277_not
g45133 not n23286 ; n23286_not
g45134 not n25194 ; n25194_not
g45135 not n23295 ; n23295_not
g45136 not n25077 ; n25077_not
g45137 not n12783 ; n12783_not
g45138 not n14790 ; n14790_not
g45139 not n12792 ; n12792_not
g45140 not n24960 ; n24960_not
g45141 not n23367 ; n23367_not
g45142 not n23394 ; n23394_not
g45143 not n14808 ; n14808_not
g45144 not n12846 ; n12846_not
g45145 not n23376 ; n23376_not
g45146 not n12828 ; n12828_not
g45147 not n23385 ; n23385_not
g45148 not n12765 ; n12765_not
g45149 not n14718 ; n14718_not
g45150 not n14835 ; n14835_not
g45151 not n25158 ; n25158_not
g45152 not n14817 ; n14817_not
g45153 not n12774 ; n12774_not
g45154 not n25149 ; n25149_not
g45155 not n14826 ; n14826_not
g45156 not n12855 ; n12855_not
g45157 not n23358 ; n23358_not
g45158 not n23349 ; n23349_not
g45159 not n14781 ; n14781_not
g45160 not n14772 ; n14772_not
g45161 not n25275 ; n25275_not
g45162 not n12936 ; n12936_not
g45163 not n15069 ; n15069_not
g45164 not n25284 ; n25284_not
g45165 not n12594 ; n12594_not
g45166 not n15078 ; n15078_not
g45167 not n12558 ; n12558_not
g45168 not n12585 ; n12585_not
g45169 not n12576 ; n12576_not
g45170 not n12945 ; n12945_not
g45171 not n15087 ; n15087_not
g45172 not n12567 ; n12567_not
g45173 not n22926 ; n22926_not
g45174 not n14709 ; n14709_not
g45175 not n12954 ; n12954_not
g45176 not n15186 ; n15186_not
g45177 not n24951 ; n24951_not
g45178 not n12972 ; n12972_not
g45179 not n25338 ; n25338_not
g45180 not n14691 ; n14691_not
g45181 not n15168 ; n15168_not
g45182 not n14682 ; n14682_not
g45183 not n23493 ; n23493_not
g45184 not n15159 ; n15159_not
g45185 not n12549 ; n12549_not
g45186 not n12963 ; n12963_not
g45187 not n14943 ; n14943_not
g45188 not n23466 ; n23466_not
g45189 not n12657 ; n12657_not
g45190 not n25248 ; n25248_not
g45191 not n25059 ; n25059_not
g45192 not n12666 ; n12666_not
g45193 not n25239 ; n25239_not
g45194 not n14925 ; n14925_not
g45195 not n14934 ; n14934_not
g45196 not n14736 ; n14736_not
g45197 not n23457 ; n23457_not
g45198 not n14916 ; n14916_not
g45199 not n23259 ; n23259_not
g45200 not n12675 ; n12675_not
g45201 not n25266 ; n25266_not
g45202 not n12918 ; n12918_not
g45203 not n23187 ; n23187_not
g45204 not n12909 ; n12909_not
g45205 not n14970 ; n14970_not
g45206 not n23178 ; n23178_not
g45207 not n12648 ; n12648_not
g45208 not n14727 ; n14727_not
g45209 not n15735 ; n15735_not
g45210 not n15744 ; n15744_not
g45211 not n24654 ; n24654_not
g45212 not n25932 ; n25932_not
g45213 not n22494 ; n22494_not
g45214 not n15753 ; n15753_not
g45215 not n22485 ; n22485_not
g45216 not n22476 ; n22476_not
g45217 not n25824 ; n25824_not
g45218 not n15762 ; n15762_not
g45219 not n14529 ; n14529_not
g45220 not n25941 ; n25941_not
g45221 not n22467 ; n22467_not
g45222 not n25950 ; n25950_not
g45223 not n11793 ; n11793_not
g45224 not n23691 ; n23691_not
g45225 not n22197 ; n22197_not
g45226 not n11829 ; n11829_not
g45227 not n15807 ; n15807_not
g45228 not n15726 ; n15726_not
g45229 not n11838 ; n11838_not
g45230 not n15780 ; n15780_not
g45231 not n25860 ; n25860_not
g45232 not n11847 ; n11847_not
g45233 not n25923 ; n25923_not
g45234 not n22458 ; n22458_not
g45235 not n15771 ; n15771_not
g45236 not n22386 ; n22386_not
g45237 not n22575 ; n22575_not
g45238 not n22566 ; n22566_not
g45239 not n24681 ; n24681_not
g45240 not n22557 ; n22557_not
g45241 not n25815 ; n25815_not
g45242 not n11883 ; n11883_not
g45243 not n22548 ; n22548_not
g45244 not n23664 ; n23664_not
g45245 not n25806 ; n25806_not
g45246 not n15708 ; n15708_not
g45247 not n22539 ; n22539_not
g45248 not n11865 ; n11865_not
g45249 not n25914 ; n25914_not
g45250 not n25851 ; n25851_not
g45251 not n23673 ; n23673_not
g45252 not n25707 ; n25707_not
g45253 not n15717 ; n15717_not
g45254 not n25770 ; n25770_not
g45255 not n24672 ; n24672_not
g45256 not n25833 ; n25833_not
g45257 not n11874 ; n11874_not
g45258 not n15870 ; n15870_not
g45259 not n22359 ; n22359_not
g45260 not n11694 ; n11694_not
g45261 not n14493 ; n14493_not
g45262 not n11676 ; n11676_not
g45263 not n11685 ; n11685_not
g45264 not n12990 ; n12990_not
g45265 not n15915 ; n15915_not
g45266 not n11667 ; n11667_not
g45267 not n15924 ; n15924_not
g45268 not n13359 ; n13359_not
g45269 not n24618 ; n24618_not
g45270 not n24609 ; n24609_not
g45271 not n22278 ; n22278_not
g45272 not n22269 ; n22269_not
g45273 not n24582 ; n24582_not
g45274 not n15582 ; n15582_not
g45275 not n23736 ; n23736_not
g45276 not n13386 ; n13386_not
g45277 not n24591 ; n24591_not
g45278 not n13377 ; n13377_not
g45279 not n22287 ; n22287_not
g45280 not n15942 ; n15942_not
g45281 not n23727 ; n23727_not
g45282 not n11595 ; n11595_not
g45283 not n14484 ; n14484_not
g45284 not n22296 ; n22296_not
g45285 not n11649 ; n11649_not
g45286 not n11748 ; n11748_not
g45287 not n15843 ; n15843_not
g45288 not n11757 ; n11757_not
g45289 not n11766 ; n11766_not
g45290 not n26058 ; n26058_not
g45291 not n24636 ; n24636_not
g45292 not n15834 ; n15834_not
g45293 not n26049 ; n26049_not
g45294 not n15825 ; n15825_not
g45295 not n11784 ; n11784_not
g45296 not n11478 ; n11478_not
g45297 not n13269 ; n13269_not
g45298 not n24627 ; n24627_not
g45299 not n26067 ; n26067_not
g45300 not n15672 ; n15672_not
g45301 not n26085 ; n26085_not
g45302 not n13287 ; n13287_not
g45303 not n22377 ; n22377_not
g45304 not n11739 ; n11739_not
g45305 not n23646 ; n23646_not
g45306 not n26076 ; n26076_not
g45307 not n22395 ; n22395_not
g45308 not n22764 ; n22764_not
g45309 not n15537 ; n15537_not
g45310 not n22755 ; n22755_not
g45311 not n25581 ; n25581_not
g45312 not n25590 ; n25590_not
g45313 not n22746 ; n22746_not
g45314 not n15546 ; n15546_not
g45315 not n14565 ; n14565_not
g45316 not n25608 ; n25608_not
g45317 not n11973 ; n11973_not
g45318 not n22737 ; n22737_not
g45319 not n13089 ; n13089_not
g45320 not n25617 ; n25617_not
g45321 not n22692 ; n22692_not
g45322 not n25653 ; n25653_not
g45323 not n23619 ; n23619_not
g45324 not n11955 ; n11955_not
g45325 not n15573 ; n15573_not
g45326 not n25644 ; n25644_not
g45327 not n25635 ; n25635_not
g45328 not n22719 ; n22719_not
g45329 not n15564 ; n15564_not
g45330 not n24726 ; n24726_not
g45331 not n24717 ; n24717_not
g45332 not n14583 ; n14583_not
g45333 not n15555 ; n15555_not
g45334 not n11964 ; n11964_not
g45335 not n11991 ; n11991_not
g45336 not n23592 ; n23592_not
g45337 not n15519 ; n15519_not
g45338 not n15492 ; n15492_not
g45339 not n22728 ; n22728_not
g45340 not n25545 ; n25545_not
g45341 not n24762 ; n24762_not
g45342 not n25536 ; n25536_not
g45343 not n22809 ; n22809_not
g45344 not n11856 ; n11856_not
g45345 not n14592 ; n14592_not
g45346 not n24771 ; n24771_not
g45347 not n15528 ; n15528_not
g45348 not n22773 ; n22773_not
g45349 not n25572 ; n25572_not
g45350 not n24744 ; n24744_not
g45351 not n11982 ; n11982_not
g45352 not n25563 ; n25563_not
g45353 not n25554 ; n25554_not
g45354 not n22791 ; n22791_not
g45355 not n24753 ; n24753_not
g45356 not n25725 ; n25725_not
g45357 not n22629 ; n22629_not
g45358 not n23637 ; n23637_not
g45359 not n15645 ; n15645_not
g45360 not n13179 ; n13179_not
g45361 not n15654 ; n15654_not
g45362 not n24708 ; n24708_not
g45363 not n25734 ; n25734_not
g45364 not n15663 ; n15663_not
g45365 not n25761 ; n25761_not
g45366 not n13197 ; n13197_not
g45367 not n14547 ; n14547_not
g45368 not n25752 ; n25752_not
g45369 not n23655 ; n23655_not
g45370 not n22593 ; n22593_not
g45371 not n13188 ; n13188_not
g45372 not n25743 ; n25743_not
g45373 not n14556 ; n14556_not
g45374 not n11919 ; n11919_not
g45375 not n22656 ; n22656_not
g45376 not n25680 ; n25680_not
g45377 not n25671 ; n25671_not
g45378 not n22647 ; n22647_not
g45379 not n15591 ; n15591_not
g45380 not n14574 ; n14574_not
g45381 not n22449 ; n22449_not
g45382 not n22665 ; n22665_not
g45383 not n22674 ; n22674_not
g45384 not n25662 ; n25662_not
g45385 not n23628 ; n23628_not
g45386 not n22683 ; n22683_not
g45387 not n25626 ; n25626_not
g45388 not n15636 ; n15636_not
g45389 not n25716 ; n25716_not
g45390 not n22638 ; n22638_not
g45391 not n11937 ; n11937_not
g45392 not n11928 ; n11928_not
g45393 not n15618 ; n15618_not
g45394 not n11892 ; n11892_not
g45395 not n15609 ; n15609_not
g45396 not n11946 ; n11946_not
g45397 not n17409 ; n17409_not
g45398 not n18174 ; n18174_not
g45399 not n17553 ; n17553_not
g45400 not n19308 ; n19308_not
g45401 not n17418 ; n17418_not
g45402 not n20775 ; n20775_not
g45403 not n19830 ; n19830_not
g45404 not n19614 ; n19614_not
g45405 not n17670 ; n17670_not
g45406 not n18381 ; n18381_not
g45407 not n17247 ; n17247_not
g45408 not n19650 ; n19650_not
g45409 not n17940 ; n17940_not
g45410 not n19506 ; n19506_not
g45411 not n20397 ; n20397_not
g45412 not n19245 ; n19245_not
g45413 not n18147 ; n18147_not
g45414 not n20757 ; n20757_not
g45415 not n18921 ; n18921_not
g45416 not n18543 ; n18543_not
g45417 not n19605 ; n19605_not
g45418 not n20874 ; n20874_not
g45419 not n19164 ; n19164_not
g45420 not n18552 ; n18552_not
g45421 not n20766 ; n20766_not
g45422 not n19371 ; n19371_not
g45423 not n18282 ; n18282_not
g45424 not n20883 ; n20883_not
g45425 not n18525 ; n18525_not
g45426 not n20838 ; n20838_not
g45427 not n19065 ; n19065_not
g45428 not n17805 ; n17805_not
g45429 not n18813 ; n18813_not
g45430 not n19155 ; n19155_not
g45431 not n20685 ; n20685_not
g45432 not n17094 ; n17094_not
g45433 not n20784 ; n20784_not
g45434 not n20658 ; n20658_not
g45435 not n21279 ; n21279_not
g45436 not n18273 ; n18273_not
g45437 not n17427 ; n17427_not
g45438 not n17256 ; n17256_not
g45439 not n17058 ; n17058_not
g45440 not n19623 ; n19623_not
g45441 not n19731 ; n19731_not
g45442 not n18471 ; n18471_not
g45443 not n19119 ; n19119_not
g45444 not n17265 ; n17265_not
g45445 not n17436 ; n17436_not
g45446 not n20649 ; n20649_not
g45447 not n17049 ; n17049_not
g45448 not n21288 ; n21288_not
g45449 not n19128 ; n19128_not
g45450 not n18336 ; n18336_not
g45451 not n17445 ; n17445_not
g45452 not n18084 ; n18084_not
g45453 not n18435 ; n18435_not
g45454 not n17841 ; n17841_not
g45455 not n20496 ; n20496_not
g45456 not n20667 ; n20667_not
g45457 not n19236 ; n19236_not
g45458 not n19146 ; n19146_not
g45459 not n17355 ; n17355_not
g45460 not n17076 ; n17076_not
g45461 not n18462 ; n18462_not
g45462 not n18129 ; n18129_not
g45463 not n19551 ; n19551_not
g45464 not n17067 ; n17067_not
g45465 not n19713 ; n19713_not
g45466 not n19137 ; n19137_not
g45467 not n18444 ; n18444_not
g45468 not n21189 ; n21189_not
g45469 not n17625 ; n17625_not
g45470 not n18291 ; n18291_not
g45471 not n19533 ; n19533_not
g45472 not n19173 ; n19173_not
g45473 not n18480 ; n18480_not
g45474 not n18831 ; n18831_not
g45475 not n18255 ; n18255_not
g45476 not n20379 ; n20379_not
g45477 not n19191 ; n19191_not
g45478 not n19740 ; n19740_not
g45479 not n18246 ; n18246_not
g45480 not n20856 ; n20856_not
g45481 not n17193 ; n17193_not
g45482 not n19263 ; n19263_not
g45483 not n18318 ; n18318_not
g45484 not n19452 ; n19452_not
g45485 not n20748 ; n20748_not
g45486 not n18183 ; n18183_not
g45487 not n18930 ; n18930_not
g45488 not n19272 ; n19272_not
g45489 not n20937 ; n20937_not
g45490 not n17373 ; n17373_not
g45491 not n17616 ; n17616_not
g45492 not n21198 ; n21198_not
g45493 not n20739 ; n20739_not
g45494 not n18327 ; n18327_not
g45495 not n18840 ; n18840_not
g45496 not n19182 ; n19182_not
g45497 not n17607 ; n17607_not
g45498 not n19524 ; n19524_not
g45499 not n17157 ; n17157_not
g45500 not n17661 ; n17661_not
g45501 not n20676 ; n20676_not
g45502 not n19542 ; n19542_not
g45503 not n17148 ; n17148_not
g45504 not n17139 ; n17139_not
g45505 not n17535 ; n17535_not
g45506 not n18057 ; n18057_not
g45507 not n18354 ; n18354_not
g45508 not n19290 ; n19290_not
g45509 not n18624 ; n18624_not
g45510 not n19254 ; n19254_not
g45511 not n19515 ; n19515_not
g45512 not n20694 ; n20694_not
g45513 not n17544 ; n17544_not
g45514 not n19902 ; n19902_not
g45515 not n17643 ; n17643_not
g45516 not n18048 ; n18048_not
g45517 not n17634 ; n17634_not
g45518 not n17184 ; n17184_not
g45519 not n19281 ; n19281_not
g45520 not n20865 ; n20865_not
g45521 not n19722 ; n19722_not
g45522 not n17760 ; n17760_not
g45523 not n17382 ; n17382_not
g45524 not n17391 ; n17391_not
g45525 not n17175 ; n17175_not
g45526 not n17166 ; n17166_not
g45527 not n17814 ; n17814_not
g45528 not n20298 ; n20298_not
g45529 not n17229 ; n17229_not
g45530 not n19218 ; n19218_not
g45531 not n19029 ; n19029_not
g45532 not n18723 ; n18723_not
g45533 not n17274 ; n17274_not
g45534 not n19083 ; n19083_not
g45535 not n20559 ; n20559_not
g45536 not n20478 ; n20478_not
g45537 not n18156 ; n18156_not
g45538 not n18642 ; n18642_not
g45539 not n19812 ; n19812_not
g45540 not n17580 ; n17580_not
g45541 not n19443 ; n19443_not
g45542 not n18417 ; n18417_not
g45543 not n19632 ; n19632_not
g45544 not n18633 ; n18633_not
g45545 not n20982 ; n20982_not
g45546 not n19047 ; n19047_not
g45547 not n20586 ; n20586_not
g45548 not n17328 ; n17328_not
g45549 not n17319 ; n17319_not
g45550 not n18237 ; n18237_not
g45551 not n18570 ; n18570_not
g45552 not n20991 ; n20991_not
g45553 not n17490 ; n17490_not
g45554 not n19092 ; n19092_not
g45555 not n20928 ; n20928_not
g45556 not n18732 ; n18732_not
g45557 not n18705 ; n18705_not
g45558 not n18426 ; n18426_not
g45559 not n20919 ; n20919_not
g45560 not n19380 ; n19380_not
g45561 not n19803 ; n19803_not
g45562 not n18309 ; n18309_not
g45563 not n17571 ; n17571_not
g45564 not n17913 ; n17913_not
g45565 not n19704 ; n19704_not
g45566 not n20568 ; n20568_not
g45567 not n19074 ; n19074_not
g45568 not n18507 ; n18507_not
g45569 not n19821 ; n19821_not
g45570 not n18165 ; n18165_not
g45571 not n19425 ; n19425_not
g45572 not n19911 ; n19911_not
g45573 not n20964 ; n20964_not
g45574 not n17472 ; n17472_not
g45575 not n20955 ; n20955_not
g45576 not n19434 ; n19434_not
g45577 not n19209 ; n19209_not
g45578 not n18903 ; n18903_not
g45579 not n19056 ; n19056_not
g45580 not n20946 ; n20946_not
g45581 not n18714 ; n18714_not
g45582 not n17283 ; n17283_not
g45583 not n18345 ; n18345_not
g45584 not n20973 ; n20973_not
g45585 not n18408 ; n18408_not
g45586 not n18912 ; n18912_not
g45587 not n18363 ; n18363_not
g45588 not n20577 ; n20577_not
g45589 not n18390 ; n18390_not
g45590 not n18264 ; n18264_not
g45591 not n18615 ; n18615_not
g45592 not n17526 ; n17526_not
g45593 not n20829 ; n20829_not
g45594 not n17454 ; n17454_not
g45595 not n17562 ; n17562_not
g45596 not n19227 ; n19227_not
g45597 not n17733 ; n17733_not
g45598 not n17517 ; n17517_not
g45599 not n17904 ; n17904_not
g45600 not n18219 ; n18219_not
g45601 not n18453 ; n18453_not
g45602 not n17742 ; n17742_not
g45603 not n18561 ; n18561_not
g45604 not n18750 ; n18750_not
g45605 not n19335 ; n19335_not
g45606 not n18534 ; n18534_not
g45607 not n18606 ; n18606_not
g45608 not n17346 ; n17346_not
g45609 not n18093 ; n18093_not
g45610 not n20892 ; n20892_not
g45611 not n17706 ; n17706_not
g45612 not n21297 ; n21297_not
g45613 not n18192 ; n18192_not
g45614 not n18651 ; n18651_not
g45615 not n19344 ; n19344_not
g45616 not n17337 ; n17337_not
g45617 not n19641 ; n19641_not
g45618 not n19353 ; n19353_not
g45619 not n20793 ; n20793_not
g45620 not n17751 ; n17751_not
g45621 not n17850 ; n17850_not
g45622 not n19461 ; n19461_not
g45623 not n19416 ; n19416_not
g45624 not n17931 ; n17931_not
g45625 not n17508 ; n17508_not
g45626 not n18066 ; n18066_not
g45627 not n18138 ; n18138_not
g45628 not n20469 ; n20469_not
g45629 not n20595 ; n20595_not
g45630 not n18228 ; n18228_not
g45631 not n19470 ; n19470_not
g45632 not n12838 ; n12838_not
g45633 not n19570 ; n19570_not
g45634 not n15844 ; n15844_not
g45635 not n22396 ; n22396_not
g45636 not n14494 ; n14494_not
g45637 not n25627 ; n25627_not
g45638 not n17572 ; n17572_not
g45639 not n12856 ; n12856_not
g45640 not n25942 ; n25942_not
g45641 not n13783 ; n13783_not
g45642 not n11866 ; n11866_not
g45643 not n25960 ; n25960_not
g45644 not n24277 ; n24277_not
g45645 not n17536 ; n17536_not
g45646 not n18256 ; n18256_not
g45647 not n24934 ; n24934_not
g45648 not n22369 ; n22369_not
g45649 not n12784 ; n12784_not
g45650 not n25906 ; n25906_not
g45651 not n15835 ; n15835_not
g45652 not n25951 ; n25951_not
g45653 not n12496 ; n12496_not
g45654 not n25915 ; n25915_not
g45655 not n14386 ; n14386_not
g45656 not n25852 ; n25852_not
g45657 not n22387 ; n22387_not
g45658 not n15817 ; n15817_not
g45659 not n25870 ; n25870_not
g45660 not n12829 ; n12829_not
g45661 not n15079 ; n15079_not
g45662 not n17509 ; n17509_not
g45663 not n17554 ; n17554_not
g45664 not n19192 ; n19192_not
g45665 not n25933 ; n25933_not
g45666 not n20839 ; n20839_not
g45667 not n15556 ; n15556_not
g45668 not n20569 ; n20569_not
g45669 not n15088 ; n15088_not
g45670 not n15808 ; n15808_not
g45671 not n25843 ; n25843_not
g45672 not n25096 ; n25096_not
g45673 not n15646 ; n15646_not
g45674 not n20848 ; n20848_not
g45675 not n13378 ; n13378_not
g45676 not n25861 ; n25861_not
g45677 not n12775 ; n12775_not
g45678 not n15826 ; n15826_not
g45679 not n23818 ; n23818_not
g45680 not n12847 ; n12847_not
g45681 not n22378 ; n22378_not
g45682 not n12793 ; n12793_not
g45683 not n15871 ; n15871_not
g45684 not n15853 ; n15853_not
g45685 not n17527 ; n17527_not
g45686 not n15862 ; n15862_not
g45687 not n16078 ; n16078_not
g45688 not n14944 ; n14944_not
g45689 not n17347 ; n17347_not
g45690 not n17518 ; n17518_not
g45691 not n16087 ; n16087_not
g45692 not n22189 ; n22189_not
g45693 not n11578 ; n11578_not
g45694 not n16096 ; n16096_not
g45695 not n17905 ; n17905_not
g45696 not n11569 ; n11569_not
g45697 not n20695 ; n20695_not
g45698 not n13828 ; n13828_not
g45699 not n11677 ; n11677_not
g45700 not n18337 ; n18337_not
g45701 not n12964 ; n12964_not
g45702 not n11668 ; n11668_not
g45703 not n19129 ; n19129_not
g45704 not n11659 ; n11659_not
g45705 not n19624 ; n19624_not
g45706 not n11596 ; n11596_not
g45707 not n18607 ; n18607_not
g45708 not n12973 ; n12973_not
g45709 not n20893 ; n20893_not
g45710 not n23692 ; n23692_not
g45711 not n23845 ; n23845_not
g45712 not n21955 ; n21955_not
g45713 not n16069 ; n16069_not
g45714 not n15691 ; n15691_not
g45715 not n22198 ; n22198_not
g45716 not n16177 ; n16177_not
g45717 not n19642 ; n19642_not
g45718 not n26176 ; n26176_not
g45719 not n14368 ; n14368_not
g45720 not n16186 ; n16186_not
g45721 not n14917 ; n14917_not
g45722 not n16195 ; n16195_not
g45723 not n19075 ; n19075_not
g45724 not n20947 ; n20947_not
g45725 not n17914 ; n17914_not
g45726 not n26194 ; n26194_not
g45727 not n24952 ; n24952_not
g45728 not n23854 ; n23854_not
g45729 not n17473 ; n17473_not
g45730 not n20956 ; n20956_not
g45731 not n16249 ; n16249_not
g45732 not n24826 ; n24826_not
g45733 not n24970 ; n24970_not
g45734 not n19093 ; n19093_not
g45735 not n26149 ; n26149_not
g45736 not n17491 ; n17491_not
g45737 not n20929 ; n20929_not
g45738 not n11497 ; n11497_not
g45739 not n26158 ; n26158_not
g45740 not n26167 ; n26167_not
g45741 not n16159 ; n16159_not
g45742 not n18238 ; n18238_not
g45743 not n19084 ; n19084_not
g45744 not n18625 ; n18625_not
g45745 not n14935 ; n14935_not
g45746 not n13189 ; n13189_not
g45747 not n16168 ; n16168_not
g45748 not n14926 ; n14926_not
g45749 not n24961 ; n24961_not
g45750 not n12883 ; n12883_not
g45751 not n15925 ; n15925_not
g45752 not n20866 ; n20866_not
g45753 not n18067 ; n18067_not
g45754 not n11794 ; n11794_not
g45755 not n18580 ; n18580_not
g45756 not n19372 ; n19372_not
g45757 not n19606 ; n19606_not
g45758 not n23188 ; n23188_not
g45759 not n11785 ; n11785_not
g45760 not n11479 ; n11479_not
g45761 not n15934 ; n15934_not
g45762 not n24097 ; n24097_not
g45763 not n22297 ; n22297_not
g45764 not n18328 ; n18328_not
g45765 not n23746 ; n23746_not
g45766 not n23827 ; n23827_not
g45767 not n25924 ; n25924_not
g45768 not n12865 ; n12865_not
g45769 not n11848 ; n11848_not
g45770 not n15880 ; n15880_not
g45771 not n13666 ; n13666_not
g45772 not n19183 ; n19183_not
g45773 not n25078 ; n25078_not
g45774 not n12874 ; n12874_not
g45775 not n15907 ; n15907_not
g45776 not n18247 ; n18247_not
g45777 not n19174 ; n19174_not
g45778 not n23179 ; n23179_not
g45779 not n15916 ; n15916_not
g45780 not n24259 ; n24259_not
g45781 not n17545 ; n17545_not
g45782 not n12937 ; n12937_not
g45783 not n26077 ; n26077_not
g45784 not n19921 ; n19921_not
g45785 not n19138 ; n19138_not
g45786 not n13639 ; n13639_not
g45787 not n19147 ; n19147_not
g45788 not n26086 ; n26086_not
g45789 not n12946 ; n12946_not
g45790 not n14962 ; n14962_not
g45791 not n18463 ; n18463_not
g45792 not n11695 ; n11695_not
g45793 not n26095 ; n26095_not
g45794 not n15970 ; n15970_not
g45795 not n12955 ; n12955_not
g45796 not n13819 ; n13819_not
g45797 not n11686 ; n11686_not
g45798 not n20875 ; n20875_not
g45799 not n11776 ; n11776_not
g45800 not n15943 ; n15943_not
g45801 not n14971 ; n14971_not
g45802 not n19165 ; n19165_not
g45803 not n13657 ; n13657_not
g45804 not n11767 ; n11767_not
g45805 not n22288 ; n22288_not
g45806 not n22279 ; n22279_not
g45807 not n12919 ; n12919_not
g45808 not n11758 ; n11758_not
g45809 not n12928 ; n12928_not
g45810 not n13765 ; n13765_not
g45811 not n26068 ; n26068_not
g45812 not n19156 ; n19156_not
g45813 not n13738 ; n13738_not
g45814 not n20884 ; n20884_not
g45815 not n11749 ; n11749_not
g45816 not n15961 ; n15961_not
g45817 not n17707 ; n17707_not
g45818 not n19048 ; n19048_not
g45819 not n18274 ; n18274_not
g45820 not n22783 ; n22783_not
g45821 not n25276 ; n25276_not
g45822 not n13387 ; n13387_not
g45823 not n11839 ; n11839_not
g45824 not n15529 ; n15529_not
g45825 not n18193 ; n18193_not
g45826 not n19336 ; n19336_not
g45827 not n18535 ; n18535_not
g45828 not n25285 ; n25285_not
g45829 not n22774 ; n22774_not
g45830 not n17680 ; n17680_not
g45831 not n19327 ; n19327_not
g45832 not n19732 ; n19732_not
g45833 not n25528 ; n25528_not
g45834 not n22765 ; n22765_not
g45835 not n19318 ; n19318_not
g45836 not n25384 ; n25384_not
g45837 not n25483 ; n25483_not
g45838 not n12199 ; n12199_not
g45839 not n17734 ; n17734_not
g45840 not n17725 ; n17725_not
g45841 not n19480 ; n19480_not
g45842 not n12577 ; n12577_not
g45843 not n15493 ; n15493_not
g45844 not n12586 ; n12586_not
g45845 not n18265 ; n18265_not
g45846 not n25492 ; n25492_not
g45847 not n22990 ; n22990_not
g45848 not n17716 ; n17716_not
g45849 not n19354 ; n19354_not
g45850 not n25294 ; n25294_not
g45851 not n23755 ; n23755_not
g45852 not n18427 ; n18427_not
g45853 not n19345 ; n19345_not
g45854 not n22792 ; n22792_not
g45855 not n19309 ; n19309_not
g45856 not n25555 ; n25555_not
g45857 not n25258 ; n25258_not
g45858 not n19507 ; n19507_not
g45859 not n15565 ; n15565_not
g45860 not n15349 ; n15349_not
g45861 not n17671 ; n17671_not
g45862 not n25474 ; n25474_not
g45863 not n12649 ; n12649_not
g45864 not n22981 ; n22981_not
g45865 not n25564 ; n25564_not
g45866 not n20686 ; n20686_not
g45867 not n11983 ; n11983_not
g45868 not n17806 ; n17806_not
g45869 not n25573 ; n25573_not
g45870 not n25582 ; n25582_not
g45871 not n18391 ; n18391_not
g45872 not n25537 ; n25537_not
g45873 not n15538 ; n15538_not
g45874 not n22756 ; n22756_not
g45875 not n20659 ; n20659_not
g45876 not n12478 ; n12478_not
g45877 not n15367 ; n15367_not
g45878 not n18490 ; n18490_not
g45879 not n14458 ; n14458_not
g45880 not n18283 ; n18283_not
g45881 not n22747 ; n22747_not
g45882 not n13729 ; n13729_not
g45883 not n15358 ; n15358_not
g45884 not n18544 ; n18544_not
g45885 not n25546 ; n25546_not
g45886 not n22738 ; n22738_not
g45887 not n20668 ; n20668_not
g45888 not n25267 ; n25267_not
g45889 not n11992 ; n11992_not
g45890 not n22729 ; n22729_not
g45891 not n22936 ; n22936_not
g45892 not n15439 ; n15439_not
g45893 not n13684 ; n13684_not
g45894 not n17761 ; n17761_not
g45895 not n12397 ; n12397_not
g45896 not n12469 ; n12469_not
g45897 not n22891 ; n22891_not
g45898 not n12379 ; n12379_not
g45899 not n19264 ; n19264_not
g45900 not n12388 ; n12388_not
g45901 not n25357 ; n25357_not
g45902 not n19390 ; n19390_not
g45903 not n22945 ; n22945_not
g45904 not n22882 ; n22882_not
g45905 not n20587 ; n20587_not
g45906 not n19444 ; n19444_not
g45907 not n19282 ; n19282_not
g45908 not n25429 ; n25429_not
g45909 not n15385 ; n15385_not
g45910 not n25375 ; n25375_not
g45911 not n14467 ; n14467_not
g45912 not n17392 ; n17392_not
g45913 not n19426 ; n19426_not
g45914 not n14476 ; n14476_not
g45915 not n22918 ; n22918_not
g45916 not n22927 ; n22927_not
g45917 not n17419 ; n17419_not
g45918 not n25393 ; n25393_not
g45919 not n19417 ; n19417_not
g45920 not n19435 ; n19435_not
g45921 not n17770 ; n17770_not
g45922 not n22909 ; n22909_not
g45923 not n24367 ; n24367_not
g45924 not n18508 ; n18508_not
g45925 not n22666 ; n22666_not
g45926 not n20578 ; n20578_not
g45927 not n19066 ; n19066_not
g45928 not n25366 ; n25366_not
g45929 not n22846 ; n22846_not
g45930 not n20596 ; n20596_not
g45931 not n22837 ; n22837_not
g45932 not n15466 ; n15466_not
g45933 not n25186 ; n25186_not
g45934 not n25339 ; n25339_not
g45935 not n12289 ; n12289_not
g45936 not n19462 ; n19462_not
g45937 not n15475 ; n15475_not
g45938 not n25465 ; n25465_not
g45939 not n22828 ; n22828_not
g45940 not n19471 ; n19471_not
g45941 not n24349 ; n24349_not
g45942 not n19363 ; n19363_not
g45943 not n24376 ; n24376_not
g45944 not n17743 ; n17743_not
g45945 not n19453 ; n19453_not
g45946 not n12568 ; n12568_not
g45947 not n22873 ; n22873_not
g45948 not n15277 ; n15277_not
g45949 not n12487 ; n12487_not
g45950 not n11947 ; n11947_not
g45951 not n11956 ; n11956_not
g45952 not n19381 ; n19381_not
g45953 not n25438 ; n25438_not
g45954 not n22864 ; n22864_not
g45955 not n25348 ; n25348_not
g45956 not n15448 ; n15448_not
g45957 not n22855 ; n22855_not
g45958 not n12298 ; n12298_not
g45959 not n15457 ; n15457_not
g45960 not n25447 ; n25447_not
g45961 not n22963 ; n22963_not
g45962 not n25195 ; n25195_not
g45963 not n23089 ; n23089_not
g45964 not n20776 ; n20776_not
g45965 not n15718 ; n15718_not
g45966 not n20497 ; n20497_not
g45967 not n19237 ; n19237_not
g45968 not n15727 ; n15727_not
g45969 not n25753 ; n25753_not
g45970 not n19552 ; n19552_not
g45971 not n12748 ; n12748_not
g45972 not n20785 ; n20785_not
g45973 not n23098 ; n23098_not
g45974 not n15745 ; n15745_not
g45975 not n19228 ; n19228_not
g45976 not n18472 ; n18472_not
g45977 not n24394 ; n24394_not
g45978 not n15736 ; n15736_not
g45979 not n15187 ; n15187_not
g45980 not n18553 ; n18553_not
g45981 not n25717 ; n25717_not
g45982 not n24268 ; n24268_not
g45983 not n11929 ; n11929_not
g45984 not n23791 ; n23791_not
g45985 not n22558 ; n22558_not
g45986 not n20758 ; n20758_not
g45987 not n25726 ; n25726_not
g45988 not n17842 ; n17842_not
g45989 not n12739 ; n12739_not
g45990 not n19255 ; n19255_not
g45991 not n11893 ; n11893_not
g45992 not n19543 ; n19543_not
g45993 not n17239 ; n17239_not
g45994 not n17590 ; n17590_not
g45995 not n20767 ; n20767_not
g45996 not n15709 ; n15709_not
g45997 not n25735 ; n25735_not
g45998 not n15169 ; n15169_not
g45999 not n25825 ; n25825_not
g46000 not n19219 ; n19219_not
g46001 not n20479 ; n20479_not
g46002 not n15772 ; n15772_not
g46003 not n19561 ; n19561_not
g46004 not n22459 ; n22459_not
g46005 not n17581 ; n17581_not
g46006 not n11875 ; n11875_not
g46007 not n12766 ; n12766_not
g46008 not n17860 ; n17860_not
g46009 not n14449 ; n14449_not
g46010 not n15781 ; n15781_not
g46011 not n12757 ; n12757_not
g46012 not n25159 ; n25159_not
g46013 not n25771 ; n25771_not
g46014 not n25780 ; n25780_not
g46015 not n22495 ; n22495_not
g46016 not n20794 ; n20794_not
g46017 not n17851 ; n17851_not
g46018 not n25672 ; n25672_not
g46019 not n13774 ; n13774_not
g46020 not n22486 ; n22486_not
g46021 not n20488 ; n20488_not
g46022 not n25807 ; n25807_not
g46023 not n15178 ; n15178_not
g46024 not n24295 ; n24295_not
g46025 not n22477 ; n22477_not
g46026 not n18562 ; n18562_not
g46027 not n22954 ; n22954_not
g46028 not n15763 ; n15763_not
g46029 not n25177 ; n25177_not
g46030 not n22468 ; n22468_not
g46031 not n18571 ; n18571_not
g46032 not n15592 ; n15592_not
g46033 not n12667 ; n12667_not
g46034 not n18481 ; n18481_not
g46035 not n11857 ; n11857_not
g46036 not n22657 ; n22657_not
g46037 not n19525 ; n19525_not
g46038 not n25636 ; n25636_not
g46039 not n15295 ; n15295_not
g46040 not n22648 ; n22648_not
g46041 not n17815 ; n17815_not
g46042 not n25645 ; n25645_not
g46043 not n13756 ; n13756_not
g46044 not n24178 ; n24178_not
g46045 not n12676 ; n12676_not
g46046 not n15286 ; n15286_not
g46047 not n17644 ; n17644_not
g46048 not n15628 ; n15628_not
g46049 not n25591 ; n25591_not
g46050 not n13747 ; n13747_not
g46051 not n23728 ; n23728_not
g46052 not n25609 ; n25609_not
g46053 not n19516 ; n19516_not
g46054 not n22684 ; n22684_not
g46055 not n11974 ; n11974_not
g46056 not n17662 ; n17662_not
g46057 not n19291 ; n19291_not
g46058 not n20677 ; n20677_not
g46059 not n15583 ; n15583_not
g46060 not n11965 ; n11965_not
g46061 not n23773 ; n23773_not
g46062 not n13675 ; n13675_not
g46063 not n25690 ; n25690_not
g46064 not n19903 ; n19903_not
g46065 not n12694 ; n12694_not
g46066 not n17833 ; n17833_not
g46067 not n22594 ; n22594_not
g46068 not n17257 ; n17257_not
g46069 not n17608 ; n17608_not
g46070 not n15673 ; n15673_not
g46071 not n22585 ; n22585_not
g46072 not n19273 ; n19273_not
g46073 not n15259 ; n15259_not
g46074 not n20749 ; n20749_not
g46075 not n15682 ; n15682_not
g46076 not n14485 ; n14485_not
g46077 not n22567 ; n22567_not
g46078 not n22576 ; n22576_not
g46079 not n25708 ; n25708_not
g46080 not n11938 ; n11938_not
g46081 not n19534 ; n19534_not
g46082 not n17824 ; n17824_not
g46083 not n17635 ; n17635_not
g46084 not n15637 ; n15637_not
g46085 not n25663 ; n25663_not
g46086 not n24385 ; n24385_not
g46087 not n17626 ; n17626_not
g46088 not n15655 ; n15655_not
g46089 not n12658 ; n12658_not
g46090 not n23782 ; n23782_not
g46091 not n15664 ; n15664_not
g46092 not n12685 ; n12685_not
g46093 not n25681 ; n25681_not
g46094 not n16690 ; n16690_not
g46095 not n21649 ; n21649_not
g46096 not n21388 ; n21388_not
g46097 not n26752 ; n26752_not
g46098 not n26671 ; n26671_not
g46099 not n23944 ; n23944_not
g46100 not n18832 ; n18832_not
g46101 not n10597 ; n10597_not
g46102 not n14278 ; n14278_not
g46103 not n14566 ; n14566_not
g46104 not n26761 ; n26761_not
g46105 not n24646 ; n24646_not
g46106 not n16708 ; n16708_not
g46107 not n16627 ; n16627_not
g46108 not n17194 ; n17194_not
g46109 not n13972 ; n13972_not
g46110 not n17923 ; n17923_not
g46111 not n16717 ; n16717_not
g46112 not n19723 ; n19723_not
g46113 not n18850 ; n18850_not
g46114 not n26716 ; n26716_not
g46115 not n14728 ; n14728_not
g46116 not n24673 ; n24673_not
g46117 not n26725 ; n26725_not
g46118 not n13567 ; n13567_not
g46119 not n13954 ; n13954_not
g46120 not n20992 ; n20992_not
g46121 not n26707 ; n26707_not
g46122 not n23467 ; n23467_not
g46123 not n13963 ; n13963_not
g46124 not n21667 ; n21667_not
g46125 not n16681 ; n16681_not
g46126 not n18184 ; n18184_not
g46127 not n21397 ; n21397_not
g46128 not n24655 ; n24655_not
g46129 not n24475 ; n24475_not
g46130 not n26743 ; n26743_not
g46131 not n14719 ; n14719_not
g46132 not n23476 ; n23476_not
g46133 not n26815 ; n26815_not
g46134 not n21595 ; n21595_not
g46135 not n18175 ; n18175_not
g46136 not n10579 ; n10579_not
g46137 not n18670 ; n18670_not
g46138 not n26824 ; n26824_not
g46139 not n13297 ; n13297_not
g46140 not n21586 ; n21586_not
g46141 not n13990 ; n13990_not
g46142 not n14683 ; n14683_not
g46143 not n16762 ; n16762_not
g46144 not n18058 ; n18058_not
g46145 not n24628 ; n24628_not
g46146 not n21577 ; n21577_not
g46147 not n18814 ; n18814_not
g46148 not n26833 ; n26833_not
g46149 not n21568 ; n21568_not
g46150 not n19741 ; n19741_not
g46151 not n23485 ; n23485_not
g46152 not n26770 ; n26770_not
g46153 not n18382 ; n18382_not
g46154 not n16726 ; n16726_not
g46155 not n18049 ; n18049_not
g46156 not n20299 ; n20299_not
g46157 not n23494 ; n23494_not
g46158 not n17176 ; n17176_not
g46159 not n16735 ; n16735_not
g46160 not n10588 ; n10588_not
g46161 not n24637 ; n24637_not
g46162 not n17167 ; n17167_not
g46163 not n13279 ; n13279_not
g46164 not n23890 ; n23890_not
g46165 not n16744 ; n16744_not
g46166 not n14692 ; n14692_not
g46167 not n17158 ; n17158_not
g46168 not n16753 ; n16753_not
g46169 not n17149 ; n17149_not
g46170 not n21775 ; n21775_not
g46171 not n26590 ; n26590_not
g46172 not n23917 ; n23917_not
g46173 not n24727 ; n24727_not
g46174 not n13099 ; n13099_not
g46175 not n18454 ; n18454_not
g46176 not n10669 ; n10669_not
g46177 not n21766 ; n21766_not
g46178 not n26509 ; n26509_not
g46179 not n24718 ; n24718_not
g46180 not n26617 ; n26617_not
g46181 not n13927 ; n13927_not
g46182 not n18364 ; n18364_not
g46183 not n26626 ; n26626_not
g46184 not n13936 ; n13936_not
g46185 not n16591 ; n16591_not
g46186 not n14764 ; n14764_not
g46187 not n21748 ; n21748_not
g46188 not n19705 ; n19705_not
g46189 not n10687 ; n10687_not
g46190 not n26635 ; n26635_not
g46191 not n17266 ; n17266_not
g46192 not n24763 ; n24763_not
g46193 not n24754 ; n24754_not
g46194 not n16573 ; n16573_not
g46195 not n26554 ; n26554_not
g46196 not n23656 ; n23656_not
g46197 not n24466 ; n24466_not
g46198 not n21793 ; n21793_not
g46199 not n17284 ; n17284_not
g46200 not n10759 ; n10759_not
g46201 not n26563 ; n26563_not
g46202 not n14782 ; n14782_not
g46203 not n24745 ; n24745_not
g46204 not n14296 ; n14296_not
g46205 not n21784 ; n21784_not
g46206 not n26464 ; n26464_not
g46207 not n26572 ; n26572_not
g46208 not n24529 ; n24529_not
g46209 not n17275 ; n17275_not
g46210 not n26473 ; n26473_not
g46211 not n14773 ; n14773_not
g46212 not n26581 ; n26581_not
g46213 not n16924 ; n16924_not
g46214 not n16654 ; n16654_not
g46215 not n26680 ; n26680_not
g46216 not n10678 ; n10678_not
g46217 not n26644 ; n26644_not
g46218 not n16663 ; n16663_not
g46219 not n14746 ; n14746_not
g46220 not n13198 ; n13198_not
g46221 not n24691 ; n24691_not
g46222 not n18373 ; n18373_not
g46223 not n21694 ; n21694_not
g46224 not n23458 ; n23458_not
g46225 not n21685 ; n21685_not
g46226 not n23935 ; n23935_not
g46227 not n23647 ; n23647_not
g46228 not n16618 ; n16618_not
g46229 not n24709 ; n24709_not
g46230 not n14755 ; n14755_not
g46231 not n19714 ; n19714_not
g46232 not n17248 ; n17248_not
g46233 not n26653 ; n26653_not
g46234 not n23449 ; n23449_not
g46235 not n14287 ; n14287_not
g46236 not n26662 ; n26662_not
g46237 not n14737 ; n14737_not
g46238 not n13945 ; n13945_not
g46239 not n23926 ; n23926_not
g46240 not n23584 ; n23584_not
g46241 not n27067 ; n27067_not
g46242 not n18742 ; n18742_not
g46243 not n14179 ; n14179_not
g46244 not n27139 ; n27139_not
g46245 not n16528 ; n16528_not
g46246 not n18733 ; n18733_not
g46247 not n27148 ; n27148_not
g46248 not n18445 ; n18445_not
g46249 not n13477 ; n13477_not
g46250 not n27157 ; n27157_not
g46251 not n23368 ; n23368_not
g46252 not n18139 ; n18139_not
g46253 not n13486 ; n13486_not
g46254 not n13792 ; n13792_not
g46255 not n27166 ; n27166_not
g46256 not n19804 ; n19804_not
g46257 not n18148 ; n18148_not
g46258 not n18157 ; n18157_not
g46259 not n27049 ; n27049_not
g46260 not n27058 ; n27058_not
g46261 not n16861 ; n16861_not
g46262 not n18751 ; n18751_not
g46263 not n18094 ; n18094_not
g46264 not n16870 ; n16870_not
g46265 not n23575 ; n23575_not
g46266 not n24547 ; n24547_not
g46267 not n13459 ; n13459_not
g46268 not n27076 ; n27076_not
g46269 not n13468 ; n13468_not
g46270 not n27085 ; n27085_not
g46271 not n16519 ; n16519_not
g46272 not n27094 ; n27094_not
g46273 not n27229 ; n27229_not
g46274 not n19822 ; n19822_not
g46275 not n16942 ; n16942_not
g46276 not n24493 ; n24493_not
g46277 not n27247 ; n27247_not
g46278 not n24484 ; n24484_not
g46279 not n27256 ; n27256_not
g46280 not n27238 ; n27238_not
g46281 not n27265 ; n27265_not
g46282 not n16951 ; n16951_not
g46283 not n18229 ; n18229_not
g46284 not n14188 ; n14188_not
g46285 not n27274 ; n27274_not
g46286 not n27283 ; n27283_not
g46287 not n14584 ; n14584_not
g46288 not n18166 ; n18166_not
g46289 not n13918 ; n13918_not
g46290 not n16906 ; n16906_not
g46291 not n14575 ; n14575_not
g46292 not n27175 ; n27175_not
g46293 not n18724 ; n18724_not
g46294 not n13495 ; n13495_not
g46295 not n27184 ; n27184_not
g46296 not n19813 ; n19813_not
g46297 not n27193 ; n27193_not
g46298 not n21379 ; n21379_not
g46299 not n14593 ; n14593_not
g46300 not n18715 ; n18715_not
g46301 not n18418 ; n18418_not
g46302 not n16933 ; n16933_not
g46303 not n13369 ; n13369_not
g46304 not n13558 ; n13558_not
g46305 not n16474 ; n16474_not
g46306 not n23962 ; n23962_not
g46307 not n24565 ; n24565_not
g46308 not n14269 ; n14269_not
g46309 not n26905 ; n26905_not
g46310 not n24592 ; n24592_not
g46311 not n17077 ; n17077_not
g46312 not n18805 ; n18805_not
g46313 not n16807 ; n16807_not
g46314 not n12991 ; n12991_not
g46315 not n23629 ; n23629_not
g46316 not n23539 ; n23539_not
g46317 not n10489 ; n10489_not
g46318 not n17068 ; n17068_not
g46319 not n14647 ; n14647_not
g46320 not n16816 ; n16816_not
g46321 not n21289 ; n21289_not
g46322 not n16771 ; n16771_not
g46323 not n14674 ; n14674_not
g46324 not n17095 ; n17095_not
g46325 not n23278 ; n23278_not
g46326 not n21559 ; n21559_not
g46327 not n26851 ; n26851_not
g46328 not n26842 ; n26842_not
g46329 not n16780 ; n16780_not
g46330 not n24619 ; n24619_not
g46331 not n14665 ; n14665_not
g46332 not n26860 ; n26860_not
g46333 not n16843 ; n16843_not
g46334 not n21298 ; n21298_not
g46335 not n14098 ; n14098_not
g46336 not n26923 ; n26923_not
g46337 not n23881 ; n23881_not
g46338 not n23980 ; n23980_not
g46339 not n21469 ; n21469_not
g46340 not n10399 ; n10399_not
g46341 not n16492 ; n16492_not
g46342 not n16852 ; n16852_not
g46343 not n13396 ; n13396_not
g46344 not n14629 ; n14629_not
g46345 not n23566 ; n23566_not
g46346 not n24556 ; n24556_not
g46347 not n24583 ; n24583_not
g46348 not n17059 ; n17059_not
g46349 not n16825 ; n16825_not
g46350 not n23548 ; n23548_not
g46351 not n26932 ; n26932_not
g46352 not n23863 ; n23863_not
g46353 not n14089 ; n14089_not
g46354 not n26941 ; n26941_not
g46355 not n18085 ; n18085_not
g46356 not n10498 ; n10498_not
g46357 not n26950 ; n26950_not
g46358 not n16834 ; n16834_not
g46359 not n21487 ; n21487_not
g46360 not n23971 ; n23971_not
g46361 not n14638 ; n14638_not
g46362 not n24574 ; n24574_not
g46363 not n24448 ; n24448_not
g46364 not n23836 ; n23836_not
g46365 not n26365 ; n26365_not
g46366 not n21964 ; n21964_not
g46367 not n14854 ; n14854_not
g46368 not n16456 ; n16456_not
g46369 not n17941 ; n17941_not
g46370 not n26374 ; n26374_not
g46371 not n10894 ; n10894_not
g46372 not n13882 ; n13882_not
g46373 not n24844 ; n24844_not
g46374 not n26392 ; n26392_not
g46375 not n14845 ; n14845_not
g46376 not n26347 ; n26347_not
g46377 not n21946 ; n21946_not
g46378 not n16465 ; n16465_not
g46379 not n24880 ; n24880_not
g46380 not n14863 ; n14863_not
g46381 not n17428 ; n17428_not
g46382 not n14872 ; n14872_not
g46383 not n26185 ; n26185_not
g46384 not n20398 ; n20398_not
g46385 not n13864 ; n13864_not
g46386 not n10957 ; n10957_not
g46387 not n24439 ; n24439_not
g46388 not n16447 ; n16447_not
g46389 not n21991 ; n21991_not
g46390 not n26329 ; n26329_not
g46391 not n10948 ; n10948_not
g46392 not n26338 ; n26338_not
g46393 not n10939 ; n10939_not
g46394 not n21982 ; n21982_not
g46395 not n24862 ; n24862_not
g46396 not n26275 ; n26275_not
g46397 not n26356 ; n26356_not
g46398 not n26428 ; n26428_not
g46399 not n24196 ; n24196_not
g46400 not n14827 ; n14827_not
g46401 not n26437 ; n26437_not
g46402 not n16483 ; n16483_not
g46403 not n21676 ; n21676_not
g46404 not n26419 ; n26419_not
g46405 not n17374 ; n17374_not
g46406 not n18940 ; n18940_not
g46407 not n23359 ; n23359_not
g46408 not n17950 ; n17950_not
g46409 not n26446 ; n26446_not
g46410 not n10768 ; n10768_not
g46411 not n24187 ; n24187_not
g46412 not n14818 ; n14818_not
g46413 not n16294 ; n16294_not
g46414 not n10885 ; n10885_not
g46415 not n19651 ; n19651_not
g46416 not n21937 ; n21937_not
g46417 not n14359 ; n14359_not
g46418 not n21928 ; n21928_not
g46419 not n18706 ; n18706_not
g46420 not n24835 ; n24835_not
g46421 not n10876 ; n10876_not
g46422 not n21919 ; n21919_not
g46423 not n21658 ; n21658_not
g46424 not n17383 ; n17383_not
g46425 not n10867 ; n10867_not
g46426 not n18634 ; n18634_not
g46427 not n20983 ; n20983_not
g46428 not n18643 ; n18643_not
g46429 not n18346 ; n18346_not
g46430 not n21829 ; n21829_not
g46431 not n16339 ; n16339_not
g46432 not n26239 ; n26239_not
g46433 not n10849 ; n10849_not
g46434 not n19633 ; n19633_not
g46435 not n16348 ; n16348_not
g46436 not n26248 ; n26248_not
g46437 not n16258 ; n16258_not
g46438 not n20965 ; n20965_not
g46439 not n11398 ; n11398_not
g46440 not n16267 ; n16267_not
g46441 not n14908 ; n14908_not
g46442 not n23683 ; n23683_not
g46443 not n23269 ; n23269_not
g46444 not n16276 ; n16276_not
g46445 not n11389 ; n11389_not
g46446 not n22099 ; n22099_not
g46447 not n24943 ; n24943_not
g46448 not n20974 ; n20974_not
g46449 not n19057 ; n19057_not
g46450 not n12982 ; n12982_not
g46451 not n24808 ; n24808_not
g46452 not n17455 ; n17455_not
g46453 not n24907 ; n24907_not
g46454 not n10984 ; n10984_not
g46455 not n26293 ; n26293_not
g46456 not n23872 ; n23872_not
g46457 not n13594 ; n13594_not
g46458 not n13855 ; n13855_not
g46459 not n10966 ; n10966_not
g46460 not n17446 ; n17446_not
g46461 not n16429 ; n16429_not
g46462 not n17437 ; n17437_not
g46463 not n16438 ; n16438_not
g46464 not n16357 ; n16357_not
g46465 not n23287 ; n23287_not
g46466 not n18319 ; n18319_not
g46467 not n16366 ; n16366_not
g46468 not n26257 ; n26257_not
g46469 not n24925 ; n24925_not
g46470 not n16375 ; n16375_not
g46471 not n13846 ; n13846_not
g46472 not n26266 ; n26266_not
g46473 not n19930 ; n19930_not
g46474 not n18436 ; n18436_not
g46475 not n17464 ; n17464_not
g46476 not n18661 ; n18661_not
g46477 not n26284 ; n26284_not
g46478 not n23296 ; n23296_not
g46479 not n16384 ; n16384_not
g46480 not n21865 ; n21865_not
g46481 not n24781 ; n24781_not
g46482 not n21838 ; n21838_not
g46483 not n26491 ; n26491_not
g46484 not n24169 ; n24169_not
g46485 not n21883 ; n21883_not
g46486 not n10777 ; n10777_not
g46487 not n26518 ; n26518_not
g46488 not n21856 ; n21856_not
g46489 not n24790 ; n24790_not
g46490 not n16564 ; n16564_not
g46491 not n14809 ; n14809_not
g46492 not n13909 ; n13909_not
g46493 not n23908 ; n23908_not
g46494 not n16555 ; n16555_not
g46495 not n10786 ; n10786_not
g46496 not n23395 ; n23395_not
g46497 not n16537 ; n16537_not
g46498 not n13576 ; n13576_not
g46499 not n24817 ; n24817_not
g46500 not n18760 ; n18760_not
g46501 not n17356 ; n17356_not
g46502 not n26527 ; n26527_not
g46503 not n14548 ; n14548_not
g46504 not n18922 ; n18922_not
g46505 not n18931 ; n18931_not
g46506 not n18904 ; n18904_not
g46507 not n18913 ; n18913_not
g46508 not n17338 ; n17338_not
g46509 not n19840 ; n19840_not
g46510 not n17329 ; n17329_not
g46511 not n19660 ; n19660_not
g46512 not n21847 ; n21847_not
g46513 not n21874 ; n21874_not
g46514 not n26536 ; n26536_not
g46515 not n20857 ; n20857_not
g46516 not n14791 ; n14791_not
g46517 not n13891 ; n13891_not
g46518 not n26383 ; n26383_not
g46519 not n24548 ; n24548_not
g46520 not n23693 ; n23693_not
g46521 not n17870 ; n17870_not
g46522 not n17906 ; n17906_not
g46523 not n19634 ; n19634_not
g46524 not n12785 ; n12785_not
g46525 not n13469 ; n13469_not
g46526 not n19472 ; n19472_not
g46527 not n24719 ; n24719_not
g46528 not n23576 ; n23576_not
g46529 not n19463 ; n19463_not
g46530 not n22955 ; n22955_not
g46531 not n19670 ; n19670_not
g46532 not n18491 ; n18491_not
g46533 not n18068 ; n18068_not
g46534 not n15179 ; n15179_not
g46535 not n24773 ; n24773_not
g46536 not n24584 ; n24584_not
g46537 not n22991 ; n22991_not
g46538 not n18095 ; n18095_not
g46539 not n22757 ; n22757_not
g46540 not n14765 ; n14765_not
g46541 not n24809 ; n24809_not
g46542 not n14945 ; n14945_not
g46543 not n14882 ; n14882_not
g46544 not n14639 ; n14639_not
g46545 not n12587 ; n12587_not
g46546 not n24566 ; n24566_not
g46547 not n24377 ; n24377_not
g46548 not n23558 ; n23558_not
g46549 not n23189 ; n23189_not
g46550 not n25295 ; n25295_not
g46551 not n12974 ; n12974_not
g46552 not n12983 ; n12983_not
g46553 not n25286 ; n25286_not
g46554 not n19553 ; n19553_not
g46555 not n18437 ; n18437_not
g46556 not n19823 ; n19823_not
g46557 not n14891 ; n14891_not
g46558 not n12794 ; n12794_not
g46559 not n24917 ; n24917_not
g46560 not n19706 ; n19706_not
g46561 not n12569 ; n12569_not
g46562 not n20489 ; n20489_not
g46563 not n17852 ; n17852_not
g46564 not n24980 ; n24980_not
g46565 not n23567 ; n23567_not
g46566 not n23297 ; n23297_not
g46567 not n13397 ; n13397_not
g46568 not n22982 ; n22982_not
g46569 not n24908 ; n24908_not
g46570 not n12578 ; n12578_not
g46571 not n18185 ; n18185_not
g46572 not n25367 ; n25367_not
g46573 not n17861 ; n17861_not
g46574 not n14594 ; n14594_not
g46575 not n13568 ; n13568_not
g46576 not n14918 ; n14918_not
g46577 not n24944 ; n24944_not
g46578 not n19436 ; n19436_not
g46579 not n24368 ; n24368_not
g46580 not n24485 ; n24485_not
g46581 not n22937 ; n22937_not
g46582 not n14783 ; n14783_not
g46583 not n14792 ; n14792_not
g46584 not n19616 ; n19616_not
g46585 not n24746 ; n24746_not
g46586 not n17924 ; n17924_not
g46587 not n15386 ; n15386_not
g46588 not n17735 ; n17735_not
g46589 not n14576 ; n14576_not
g46590 not n14927 ; n14927_not
g46591 not n19814 ; n19814_not
g46592 not n24953 ; n24953_not
g46593 not n25376 ; n25376_not
g46594 not n22928 ; n22928_not
g46595 not n14909 ; n14909_not
g46596 not n18167 ; n18167_not
g46597 not n18257 ; n18257_not
g46598 not n14666 ; n14666_not
g46599 not n14549 ; n14549_not
g46600 not n14585 ; n14585_not
g46601 not n18248 ; n18248_not
g46602 not n17915 ; n17915_not
g46603 not n23684 ; n23684_not
g46604 not n14729 ; n14729_not
g46605 not n24494 ; n24494_not
g46606 not n12767 ; n12767_not
g46607 not n18158 ; n18158_not
g46608 not n22856 ; n22856_not
g46609 not n24755 ; n24755_not
g46610 not n12758 ; n12758_not
g46611 not n24728 ; n24728_not
g46612 not n13667 ; n13667_not
g46613 not n14774 ; n14774_not
g46614 not n23585 ; n23585_not
g46615 not n12497 ; n12497_not
g46616 not n17780 ; n17780_not
g46617 not n14936 ; n14936_not
g46618 not n25178 ; n25178_not
g46619 not n24926 ; n24926_not
g46620 not n23288 ; n23288_not
g46621 not n22964 ; n22964_not
g46622 not n19454 ; n19454_not
g46623 not n24971 ; n24971_not
g46624 not n23387 ; n23387_not
g46625 not n19940 ; n19940_not
g46626 not n12479 ; n12479_not
g46627 not n24395 ; n24395_not
g46628 not n22946 ; n22946_not
g46629 not n23396 ; n23396_not
g46630 not n15098 ; n15098_not
g46631 not n24737 ; n24737_not
g46632 not n19427 ; n19427_not
g46633 not n13496 ; n13496_not
g46634 not n13595 ; n13595_not
g46635 not n18176 ; n18176_not
g46636 not n25169 ; n25169_not
g46637 not n23279 ; n23279_not
g46638 not n19805 ; n19805_not
g46639 not n15089 ; n15089_not
g46640 not n24764 ; n24764_not
g46641 not n13487 ; n13487_not
g46642 not n25349 ; n25349_not
g46643 not n24296 ; n24296_not
g46644 not n24962 ; n24962_not
g46645 not n15296 ; n15296_not
g46646 not n24692 ; n24692_not
g46647 not n14837 ; n14837_not
g46648 not n23495 ; n23495_not
g46649 not n24638 ; n24638_not
g46650 not n18239 ; n18239_not
g46651 not n12893 ; n12893_not
g46652 not n17816 ; n17816_not
g46653 not n14738 ; n14738_not
g46654 not n19526 ; n19526_not
g46655 not n12857 ; n12857_not
g46656 not n12884 ; n12884_not
g46657 not n14693 ; n14693_not
g46658 not n19571 ; n19571_not
g46659 not n12677 ; n12677_not
g46660 not n24836 ; n24836_not
g46661 not n24467 ; n24467_not
g46662 not n24476 ; n24476_not
g46663 not n14495 ; n14495_not
g46664 not n19742 ; n19742_not
g46665 not n23666 ; n23666_not
g46666 not n17825 ; n17825_not
g46667 not n13676 ; n13676_not
g46668 not n24845 ; n24845_not
g46669 not n23369 ; n23369_not
g46670 not n18482 ; n18482_not
g46671 not n15287 ; n15287_not
g46672 not n14846 ; n14846_not
g46673 not n13298 ; n13298_not
g46674 not n14747 ; n14747_not
g46675 not n12848 ; n12848_not
g46676 not n14972 ; n14972_not
g46677 not n17708 ; n17708_not
g46678 not n19751 ; n19751_not
g46679 not n19652 ; n19652_not
g46680 not n20498 ; n20498_not
g46681 not n19355 ; n19355_not
g46682 not n13658 ; n13658_not
g46683 not n13199 ; n13199_not
g46684 not n12992 ; n12992_not
g46685 not n19508 ; n19508_not
g46686 not n12686 ; n12686_not
g46687 not n17771 ; n17771_not
g46688 not n24386 ; n24386_not
g46689 not n19733 ; n19733_not
g46690 not n25079 ; n25079_not
g46691 not n14990 ; n14990_not
g46692 not n12866 ; n12866_not
g46693 not n24656 ; n24656_not
g46694 not n12695 ; n12695_not
g46695 not n17951 ; n17951_not
g46696 not n17834 ; n17834_not
g46697 not n24665 ; n24665_not
g46698 not n17663 ; n17663_not
g46699 not n23468 ; n23468_not
g46700 not n24629 ; n24629_not
g46701 not n14819 ; n14819_not
g46702 not n23657 ; n23657_not
g46703 not n14486 ; n14486_not
g46704 not n23486 ; n23486_not
g46705 not n12659 ; n12659_not
g46706 not n19175 ; n19175_not
g46707 not n23459 ; n23459_not
g46708 not n14828 ; n14828_not
g46709 not n25097 ; n25097_not
g46710 not n15278 ; n15278_not
g46711 not n24647 ; n24647_not
g46712 not n14567 ; n14567_not
g46713 not n12875 ; n12875_not
g46714 not n19535 ; n19535_not
g46715 not n24818 ; n24818_not
g46716 not n13577 ; n13577_not
g46717 not n24827 ; n24827_not
g46718 not n24674 ; n24674_not
g46719 not n23477 ; n23477_not
g46720 not n18446 ; n18446_not
g46721 not n12956 ; n12956_not
g46722 not n24791 ; n24791_not
g46723 not n20399 ; n20399_not
g46724 not n18194 ; n18194_not
g46725 not n12398 ; n12398_not
g46726 not n15359 ; n15359_not
g46727 not n14648 ; n14648_not
g46728 not n15188 ; n15188_not
g46729 not n19580 ; n19580_not
g46730 not n24872 ; n24872_not
g46731 not n14756 ; n14756_not
g46732 not n13559 ; n13559_not
g46733 not n18077 ; n18077_not
g46734 not n14864 ; n14864_not
g46735 not n13586 ; n13586_not
g46736 not n14963 ; n14963_not
g46737 not n24593 ; n24593_not
g46738 not n13379 ; n13379_not
g46739 not n24575 ; n24575_not
g46740 not n23729 ; n23729_not
g46741 not n14954 ; n14954_not
g46742 not n13388 ; n13388_not
g46743 not n18086 ; n18086_not
g46744 not n18473 ; n18473_not
g46745 not n12749 ; n12749_not
g46746 not n24881 ; n24881_not
g46747 not n25277 ; n25277_not
g46748 not n23099 ; n23099_not
g46749 not n19625 ; n19625_not
g46750 not n23549 ; n23549_not
g46751 not n14981 ; n14981_not
g46752 not n19643 ; n19643_not
g46753 not n19490 ; n19490_not
g46754 not n12965 ; n12965_not
g46755 not n14873 ; n14873_not
g46756 not n17807 ; n17807_not
g46757 not n14675 ; n14675_not
g46758 not n25196 ; n25196_not
g46759 not n18464 ; n18464_not
g46760 not n12839 ; n12839_not
g46761 not n13649 ; n13649_not
g46762 not n17960 ; n17960_not
g46763 not n17942 ; n17942_not
g46764 not n23198 ; n23198_not
g46765 not n15197 ; n15197_not
g46766 not n18059 ; n18059_not
g46767 not n14684 ; n14684_not
g46768 not n19517 ; n19517_not
g46769 not n23648 ; n23648_not
g46770 not n23378 ; n23378_not
g46771 not n19715 ; n19715_not
g46772 not n25259 ; n25259_not
g46773 not n24863 ; n24863_not
g46774 not n17843 ; n17843_not
g46775 not n19760 ; n19760_not
g46776 not n12938 ; n12938_not
g46777 not n24458 ; n24458_not
g46778 not n19841 ; n19841_not
g46779 not n24854 ; n24854_not
g46780 not n14855 ; n14855_not
g46781 not n24449 ; n24449_not
g46782 not n12929 ; n12929_not
g46783 not n21875 ; n21875_not
g46784 not n26492 ; n26492_not
g46785 not n21866 ; n21866_not
g46786 not n15782 ; n15782_not
g46787 not n17357 ; n17357_not
g46788 not n18914 ; n18914_not
g46789 not n21857 ; n21857_not
g46790 not n17348 ; n17348_not
g46791 not n21848 ; n21848_not
g46792 not n16529 ; n16529_not
g46793 not n21839 ; n21839_not
g46794 not n16538 ; n16538_not
g46795 not n13919 ; n13919_not
g46796 not n10787 ; n10787_not
g46797 not n16547 ; n16547_not
g46798 not n26519 ; n26519_not
g46799 not n16556 ; n16556_not
g46800 not n10778 ; n10778_not
g46801 not n26528 ; n26528_not
g46802 not n18905 ; n18905_not
g46803 not n18950 ; n18950_not
g46804 not n17384 ; n17384_not
g46805 not n26429 ; n26429_not
g46806 not n10868 ; n10868_not
g46807 not n16484 ; n16484_not
g46808 not n26438 ; n26438_not
g46809 not n18941 ; n18941_not
g46810 not n10859 ; n10859_not
g46811 not n16493 ; n16493_not
g46812 not n18932 ; n18932_not
g46813 not n26456 ; n26456_not
g46814 not n23972 ; n23972_not
g46815 not n13892 ; n13892_not
g46816 not n21893 ; n21893_not
g46817 not n26465 ; n26465_not
g46818 not n21884 ; n21884_not
g46819 not n24179 ; n24179_not
g46820 not n17366 ; n17366_not
g46821 not n26474 ; n26474_not
g46822 not n18923 ; n18923_not
g46823 not n26618 ; n26618_not
g46824 not n10697 ; n10697_not
g46825 not n13928 ; n13928_not
g46826 not n21758 ; n21758_not
g46827 not n26627 ; n26627_not
g46828 not n16592 ; n16592_not
g46829 not n21749 ; n21749_not
g46830 not n14288 ; n14288_not
g46831 not n10688 ; n10688_not
g46832 not n17267 ; n17267_not
g46833 not n18365 ; n18365_not
g46834 not n16619 ; n16619_not
g46835 not n26636 ; n26636_not
g46836 not n17258 ; n17258_not
g46837 not n13937 ; n13937_not
g46838 not n26591 ; n26591_not
g46839 not n18860 ; n18860_not
g46840 not n26645 ; n26645_not
g46841 not n17249 ; n17249_not
g46842 not n26654 ; n26654_not
g46843 not n16637 ; n16637_not
g46844 not n17294 ; n17294_not
g46845 not n26537 ; n26537_not
g46846 not n23909 ; n23909_not
g46847 not n10769 ; n10769_not
g46848 not n26555 ; n26555_not
g46849 not n21794 ; n21794_not
g46850 not n17285 ; n17285_not
g46851 not n16574 ; n16574_not
g46852 not n26564 ; n26564_not
g46853 not n14297 ; n14297_not
g46854 not n21785 ; n21785_not
g46855 not n26573 ; n26573_not
g46856 not n17276 ; n17276_not
g46857 not n26582 ; n26582_not
g46858 not n23918 ; n23918_not
g46859 not n21776 ; n21776_not
g46860 not n26609 ; n26609_not
g46861 not n18761 ; n18761_not
g46862 not n21767 ; n21767_not
g46863 not n20984 ; n20984_not
g46864 not n18644 ; n18644_not
g46865 not n18635 ; n18635_not
g46866 not n16349 ; n16349_not
g46867 not n16358 ; n16358_not
g46868 not n26249 ; n26249_not
g46869 not n18653 ; n18653_not
g46870 not n23864 ; n23864_not
g46871 not n15926 ; n15926_not
g46872 not n16367 ; n16367_not
g46873 not n17465 ; n17465_not
g46874 not n16376 ; n16376_not
g46875 not n26258 ; n26258_not
g46876 not n26276 ; n26276_not
g46877 not n17456 ; n17456_not
g46878 not n16385 ; n16385_not
g46879 not n26285 ; n26285_not
g46880 not n10985 ; n10985_not
g46881 not n16394 ; n16394_not
g46882 not n16196 ; n16196_not
g46883 not n19076 ; n19076_not
g46884 not n26186 ; n26186_not
g46885 not n20948 ; n20948_not
g46886 not n26195 ; n26195_not
g46887 not n16079 ; n16079_not
g46888 not n17474 ; n17474_not
g46889 not n23855 ; n23855_not
g46890 not n16259 ; n16259_not
g46891 not n16268 ; n16268_not
g46892 not n20966 ; n20966_not
g46893 not n11399 ; n11399_not
g46894 not n16277 ; n16277_not
g46895 not n13847 ; n13847_not
g46896 not n20957 ; n20957_not
g46897 not n20975 ; n20975_not
g46898 not n19058 ; n19058_not
g46899 not n16295 ; n16295_not
g46900 not n18347 ; n18347_not
g46901 not n23882 ; n23882_not
g46902 not n26366 ; n26366_not
g46903 not n21965 ; n21965_not
g46904 not n21956 ; n21956_not
g46905 not n26375 ; n26375_not
g46906 not n10895 ; n10895_not
g46907 not n16457 ; n16457_not
g46908 not n26384 ; n26384_not
g46909 not n26393 ; n26393_not
g46910 not n24188 ; n24188_not
g46911 not n17393 ; n17393_not
g46912 not n16466 ; n16466_not
g46913 not n21938 ; n21938_not
g46914 not n10886 ; n10886_not
g46915 not n10877 ; n10877_not
g46916 not n21929 ; n21929_not
g46917 not n16475 ; n16475_not
g46918 not n24197 ; n24197_not
g46919 not n26294 ; n26294_not
g46920 not n23873 ; n23873_not
g46921 not n10976 ; n10976_not
g46922 not n10967 ; n10967_not
g46923 not n17447 ; n17447_not
g46924 not n17438 ; n17438_not
g46925 not n16439 ; n16439_not
g46926 not n21983 ; n21983_not
g46927 not n13865 ; n13865_not
g46928 not n17429 ; n17429_not
g46929 not n16448 ; n16448_not
g46930 not n10958 ; n10958_not
g46931 not n10949 ; n10949_not
g46932 not n21992 ; n21992_not
g46933 not n26339 ; n26339_not
g46934 not n26348 ; n26348_not
g46935 not n13874 ; n13874_not
g46936 not n14099 ; n14099_not
g46937 not n26960 ; n26960_not
g46938 not n26924 ; n26924_not
g46939 not n21479 ; n21479_not
g46940 not n21299 ; n21299_not
g46941 not n26942 ; n26942_not
g46942 not n23981 ; n23981_not
g46943 not n16853 ; n16853_not
g46944 not n18770 ; n18770_not
g46945 not n18527 ; n18527_not
g46946 not n18545 ; n18545_not
g46947 not n16862 ; n16862_not
g46948 not n27059 ; n27059_not
g46949 not n16871 ; n16871_not
g46950 not n27068 ; n27068_not
g46951 not n19913 ; n19913_not
g46952 not n18806 ; n18806_not
g46953 not n26906 ; n26906_not
g46954 not n17078 ; n17078_not
g46955 not n16808 ; n16808_not
g46956 not n26915 ; n26915_not
g46957 not n17069 ; n17069_not
g46958 not n10499 ; n10499_not
g46959 not n23756 ; n23756_not
g46960 not n16826 ; n16826_not
g46961 not n16817 ; n16817_not
g46962 not n26933 ; n26933_not
g46963 not n26762 ; n26762_not
g46964 not n16736 ; n16736_not
g46965 not n26951 ; n26951_not
g46966 not n21488 ; n21488_not
g46967 not n16835 ; n16835_not
g46968 not n27176 ; n27176_not
g46969 not n16916 ; n16916_not
g46970 not n27185 ; n27185_not
g46971 not n27194 ; n27194_not
g46972 not n14189 ; n14189_not
g46973 not n16925 ; n16925_not
g46974 not n18716 ; n18716_not
g46975 not n18419 ; n18419_not
g46976 not n16934 ; n16934_not
g46977 not n18707 ; n18707_not
g46978 not n27239 ; n27239_not
g46979 not n16943 ; n16943_not
g46980 not n27248 ; n27248_not
g46981 not n18608 ; n18608_not
g46982 not n27257 ; n27257_not
g46983 not n16952 ; n16952_not
g46984 not n27275 ; n27275_not
g46985 not n16961 ; n16961_not
g46986 not n13964 ; n13964_not
g46987 not n27293 ; n27293_not
g46988 not n13856 ; n13856_not
g46989 not n27077 ; n27077_not
g46990 not n18743 ; n18743_not
g46991 not n27086 ; n27086_not
g46992 not n23963 ; n23963_not
g46993 not n16880 ; n16880_not
g46994 not n18734 ; n18734_not
g46995 not n27149 ; n27149_not
g46996 not n27158 ; n27158_not
g46997 not n23990 ; n23990_not
g46998 not n27167 ; n27167_not
g46999 not n21398 ; n21398_not
g47000 not n21389 ; n21389_not
g47001 not n18725 ; n18725_not
g47002 not n16907 ; n16907_not
g47003 not n21668 ; n21668_not
g47004 not n10598 ; n10598_not
g47005 not n16682 ; n16682_not
g47006 not n26735 ; n26735_not
g47007 not n21659 ; n21659_not
g47008 not n18374 ; n18374_not
g47009 not n26744 ; n26744_not
g47010 not n18833 ; n18833_not
g47011 not n26753 ; n26753_not
g47012 not n16691 ; n16691_not
g47013 not n16628 ; n16628_not
g47014 not n16781 ; n16781_not
g47015 not n17195 ; n17195_not
g47016 not n16709 ; n16709_not
g47017 not n20894 ; n20894_not
g47018 not n23945 ; n23945_not
g47019 not n26663 ; n26663_not
g47020 not n26672 ; n26672_not
g47021 not n26681 ; n26681_not
g47022 not n26690 ; n26690_not
g47023 not n16664 ; n16664_not
g47024 not n23927 ; n23927_not
g47025 not n21695 ; n21695_not
g47026 not n16655 ; n16655_not
g47027 not n10679 ; n10679_not
g47028 not n26708 ; n26708_not
g47029 not n21686 ; n21686_not
g47030 not n23936 ; n23936_not
g47031 not n13946 ; n13946_not
g47032 not n21677 ; n21677_not
g47033 not n18851 ; n18851_not
g47034 not n26717 ; n26717_not
g47035 not n18842 ; n18842_not
g47036 not n16673 ; n16673_not
g47037 not n26726 ; n26726_not
g47038 not n21578 ; n21578_not
g47039 not n26834 ; n26834_not
g47040 not n21569 ; n21569_not
g47041 not n17096 ; n17096_not
g47042 not n16772 ; n16772_not
g47043 not n26825 ; n26825_not
g47044 not n13991 ; n13991_not
g47045 not n26843 ; n26843_not
g47046 not n18671 ; n18671_not
g47047 not n26852 ; n26852_not
g47048 not n24089 ; n24089_not
g47049 not n18383 ; n18383_not
g47050 not n26861 ; n26861_not
g47051 not n17087 ; n17087_not
g47052 not n16790 ; n16790_not
g47053 not n26870 ; n26870_not
g47054 not n13973 ; n13973_not
g47055 not n26771 ; n26771_not
g47056 not n26780 ; n26780_not
g47057 not n16718 ; n16718_not
g47058 not n14279 ; n14279_not
g47059 not n16727 ; n16727_not
g47060 not n26807 ; n26807_not
g47061 not n17177 ; n17177_not
g47062 not n23954 ; n23954_not
g47063 not n16745 ; n16745_not
g47064 not n18824 ; n18824_not
g47065 not n17159 ; n17159_not
g47066 not n16754 ; n16754_not
g47067 not n21596 ; n21596_not
g47068 not n24098 ; n24098_not
g47069 not n21587 ; n21587_not
g47070 not n26816 ; n26816_not
g47071 not n16763 ; n16763_not
g47072 not n18815 ; n18815_not
g47073 not n22577 ; n22577_not
g47074 not n25709 ; n25709_not
g47075 not n22568 ; n22568_not
g47076 not n25718 ; n25718_not
g47077 not n19904 ; n19904_not
g47078 not n18293 ; n18293_not
g47079 not n22559 ; n22559_not
g47080 not n20759 ; n20759_not
g47081 not n15692 ; n15692_not
g47082 not n25727 ; n25727_not
g47083 not n19256 ; n19256_not
g47084 not n20597 ; n20597_not
g47085 not n19247 ; n19247_not
g47086 not n25448 ; n25448_not
g47087 not n17591 ; n17591_not
g47088 not n23792 ; n23792_not
g47089 not n25592 ; n25592_not
g47090 not n25736 ; n25736_not
g47091 not n24269 ; n24269_not
g47092 not n19229 ; n19229_not
g47093 not n25664 ; n25664_not
g47094 not n13757 ; n13757_not
g47095 not n17627 ; n17627_not
g47096 not n15647 ; n15647_not
g47097 not n15656 ; n15656_not
g47098 not n17618 ; n17618_not
g47099 not n15665 ; n15665_not
g47100 not n19274 ; n19274_not
g47101 not n25682 ; n25682_not
g47102 not n13694 ; n13694_not
g47103 not n25691 ; n25691_not
g47104 not n25457 ; n25457_not
g47105 not n22595 ; n22595_not
g47106 not n11948 ; n11948_not
g47107 not n15674 ; n15674_not
g47108 not n22586 ; n22586_not
g47109 not n11939 ; n11939_not
g47110 not n15683 ; n15683_not
g47111 not n22487 ; n22487_not
g47112 not n20795 ; n20795_not
g47113 not n25808 ; n25808_not
g47114 not n22478 ; n22478_not
g47115 not n13775 ; n13775_not
g47116 not n15377 ; n15377_not
g47117 not n24359 ; n24359_not
g47118 not n11876 ; n11876_not
g47119 not n15764 ; n15764_not
g47120 not n19373 ; n19373_not
g47121 not n12299 ; n12299_not
g47122 not n15773 ; n15773_not
g47123 not n17582 ; n17582_not
g47124 not n18572 ; n18572_not
g47125 not n25835 ; n25835_not
g47126 not n24287 ; n24287_not
g47127 not n15719 ; n15719_not
g47128 not n20777 ; n20777_not
g47129 not n13766 ; n13766_not
g47130 not n22847 ; n22847_not
g47131 not n19238 ; n19238_not
g47132 not n15728 ; n15728_not
g47133 not n25754 ; n25754_not
g47134 not n20786 ; n20786_not
g47135 not n15746 ; n15746_not
g47136 not n15737 ; n15737_not
g47137 not n11894 ; n11894_not
g47138 not n25772 ; n25772_not
g47139 not n22496 ; n22496_not
g47140 not n15755 ; n15755_not
g47141 not n25790 ; n25790_not
g47142 not n22775 ; n22775_not
g47143 not n19364 ; n19364_not
g47144 not n17690 ; n17690_not
g47145 not n19328 ; n19328_not
g47146 not n25529 ; n25529_not
g47147 not n19319 ; n19319_not
g47148 not n22766 ; n22766_not
g47149 not n15476 ; n15476_not
g47150 not n25538 ; n25538_not
g47151 not n17681 ; n17681_not
g47152 not n15539 ; n15539_not
g47153 not n22748 ; n22748_not
g47154 not n11984 ; n11984_not
g47155 not n11993 ; n11993_not
g47156 not n15557 ; n15557_not
g47157 not n25556 ; n25556_not
g47158 not n25475 ; n25475_not
g47159 not n15485 ; n15485_not
g47160 not n25484 ; n25484_not
g47161 not n17726 ; n17726_not
g47162 not n11768 ; n11768_not
g47163 not n15494 ; n15494_not
g47164 not n17744 ; n17744_not
g47165 not n22739 ; n22739_not
g47166 not n17717 ; n17717_not
g47167 not n25493 ; n25493_not
g47168 not n19346 ; n19346_not
g47169 not n22793 ; n22793_not
g47170 not n22784 ; n22784_not
g47171 not n19337 ; n19337_not
g47172 not n14459 ; n14459_not
g47173 not n18536 ; n18536_not
g47174 not n23774 ; n23774_not
g47175 not n13748 ; n13748_not
g47176 not n22658 ; n22658_not
g47177 not n17564 ; n17564_not
g47178 not n19283 ; n19283_not
g47179 not n11957 ; n11957_not
g47180 not n22649 ; n22649_not
g47181 not n15467 ; n15467_not
g47182 not n25646 ; n25646_not
g47183 not n25637 ; n25637_not
g47184 not n17654 ; n17654_not
g47185 not n14468 ; n14468_not
g47186 not n25628 ; n25628_not
g47187 not n19265 ; n19265_not
g47188 not n17645 ; n17645_not
g47189 not n15629 ; n15629_not
g47190 not n25655 ; n25655_not
g47191 not n17636 ; n17636_not
g47192 not n20678 ; n20678_not
g47193 not n15566 ; n15566_not
g47194 not n17672 ; n17672_not
g47195 not n18392 ; n18392_not
g47196 not n25565 ; n25565_not
g47197 not n23765 ; n23765_not
g47198 not n25583 ; n25583_not
g47199 not n13739 ; n13739_not
g47200 not n11966 ; n11966_not
g47201 not n11975 ; n11975_not
g47202 not n22685 ; n22685_not
g47203 not n25466 ; n25466_not
g47204 not n22676 ; n22676_not
g47205 not n20696 ; n20696_not
g47206 not n15584 ; n15584_not
g47207 not n22829 ; n22829_not
g47208 not n19049 ; n19049_not
g47209 not n22667 ; n22667_not
g47210 not n11759 ; n11759_not
g47211 not n17528 ; n17528_not
g47212 not n15953 ; n15953_not
g47213 not n26069 ; n26069_not
g47214 not n20885 ; n20885_not
g47215 not n19418 ; n19418_not
g47216 not n25385 ; n25385_not
g47217 not n15962 ; n15962_not
g47218 not n18581 ; n18581_not
g47219 not n18275 ; n18275_not
g47220 not n23837 ; n23837_not
g47221 not n19148 ; n19148_not
g47222 not n25394 ; n25394_not
g47223 not n26087 ; n26087_not
g47224 not n15971 ; n15971_not
g47225 not n19139 ; n19139_not
g47226 not n11696 ; n11696_not
g47227 not n22919 ; n22919_not
g47228 not n15980 ; n15980_not
g47229 not n22289 ; n22289_not
g47230 not n18563 ; n18563_not
g47231 not n20867 ; n20867_not
g47232 not n18428 ; n18428_not
g47233 not n19409 ; n19409_not
g47234 not n11786 ; n11786_not
g47235 not n15935 ; n15935_not
g47236 not n18266 ; n18266_not
g47237 not n13793 ; n13793_not
g47238 not n18518 ; n18518_not
g47239 not n11777 ; n11777_not
g47240 not n19166 ; n19166_not
g47241 not n22298 ; n22298_not
g47242 not n15944 ; n15944_not
g47243 not n18329 ; n18329_not
g47244 not n20876 ; n20876_not
g47245 not n18509 ; n18509_not
g47246 not n20579 ; n20579_not
g47247 not n23846 ; n23846_not
g47248 not n17519 ; n17519_not
g47249 not n16097 ; n16097_not
g47250 not n13829 ; n13829_not
g47251 not n19094 ; n19094_not
g47252 not n16088 ; n16088_not
g47253 not n17492 ; n17492_not
g47254 not n14477 ; n14477_not
g47255 not n26159 ; n26159_not
g47256 not n11498 ; n11498_not
g47257 not n26177 ; n26177_not
g47258 not n16169 ; n16169_not
g47259 not n17483 ; n17483_not
g47260 not n20939 ; n20939_not
g47261 not n18626 ; n18626_not
g47262 not n16187 ; n16187_not
g47263 not n26096 ; n26096_not
g47264 not n19922 ; n19922_not
g47265 not n11687 ; n11687_not
g47266 not n14378 ; n14378_not
g47267 not n11678 ; n11678_not
g47268 not n18338 ; n18338_not
g47269 not n11669 ; n11669_not
g47270 not n18590 ; n18590_not
g47271 not n11597 ; n11597_not
g47272 not n15863 ; n15863_not
g47273 not n14369 ; n14369_not
g47274 not n11588 ; n11588_not
g47275 not n22199 ; n22199_not
g47276 not n11579 ; n11579_not
g47277 not n25880 ; n25880_not
g47278 not n15449 ; n15449_not
g47279 not n25745 ; n25745_not
g47280 not n15845 ; n15845_not
g47281 not n11867 ; n11867_not
g47282 not n25907 ; n25907_not
g47283 not n22397 ; n22397_not
g47284 not n19382 ; n19382_not
g47285 not n22874 ; n22874_not
g47286 not n17555 ; n17555_not
g47287 not n22388 ; n22388_not
g47288 not n15854 ; n15854_not
g47289 not n22883 ; n22883_not
g47290 not n24278 ; n24278_not
g47291 not n25844 ; n25844_not
g47292 not n15791 ; n15791_not
g47293 not n25781 ; n25781_not
g47294 not n23594 ; n23594_not
g47295 not n25439 ; n25439_not
g47296 not n19067 ; n19067_not
g47297 not n15809 ; n15809_not
g47298 not n25862 ; n25862_not
g47299 not n25871 ; n25871_not
g47300 not n22865 ; n22865_not
g47301 not n15818 ; n15818_not
g47302 not n15827 ; n15827_not
g47303 not n14387 ; n14387_not
g47304 not n25952 ; n25952_not
g47305 not n25961 ; n25961_not
g47306 not n15881 ; n15881_not
g47307 not n23828 ; n23828_not
g47308 not n11849 ; n11849_not
g47309 not n15890 ; n15890_not
g47310 not n17762 ; n17762_not
g47311 not n19184 ; n19184_not
g47312 not n17537 ; n17537_not
g47313 not n15908 ; n15908_not
g47314 not n11795 ; n11795_not
g47315 not n17546 ; n17546_not
g47316 not n15917 ; n15917_not
g47317 not n20858 ; n20858_not
g47318 not n23819 ; n23819_not
g47319 not n22379 ; n22379_not
g47320 not n25925 ; n25925_not
g47321 not n11858 ; n11858_not
g47322 not n19193 ; n19193_not
g47323 not n20849 ; n20849_not
g47324 not n25934 ; n25934_not
g47325 not n13784 ; n13784_not
g47326 not n12389 ; n12389_not
g47327 not n19391 ; n19391_not
g47328 not n14199 ; n14199_not
g47329 not n17385 ; n17385_not
g47330 not n13857 ; n13857_not
g47331 not n13488 ; n13488_not
g47332 not n13938 ; n13938_not
g47333 not n13695 ; n13695_not
g47334 not n13686 ; n13686_not
g47335 not n18069 ; n18069_not
g47336 not n18429 ; n18429_not
g47337 not n23991 ; n23991_not
g47338 not n13875 ; n13875_not
g47339 not n13659 ; n13659_not
g47340 not n13758 ; n13758_not
g47341 not n24198 ; n24198_not
g47342 not n13578 ; n13578_not
g47343 not n13668 ; n13668_not
g47344 not n19932 ; n19932_not
g47345 not n13785 ; n13785_not
g47346 not n24189 ; n24189_not
g47347 not n13893 ; n13893_not
g47348 not n19950 ; n19950_not
g47349 not n24459 ; n24459_not
g47350 not n19914 ; n19914_not
g47351 not n23946 ; n23946_not
g47352 not n13596 ; n13596_not
g47353 not n13839 ; n13839_not
g47354 not n13848 ; n13848_not
g47355 not n19860 ; n19860_not
g47356 not n19851 ; n19851_not
g47357 not n24279 ; n24279_not
g47358 not n13587 ; n13587_not
g47359 not n13794 ; n13794_not
g47360 not n13866 ; n13866_not
g47361 not n19842 ; n19842_not
g47362 not n19833 ; n19833_not
g47363 not n13965 ; n13965_not
g47364 not n13974 ; n13974_not
g47365 not n13983 ; n13983_not
g47366 not n18438 ; n18438_not
g47367 not n13749 ; n13749_not
g47368 not n13992 ; n13992_not
g47369 not n19824 ; n19824_not
g47370 not n24378 ; n24378_not
g47371 not n13398 ; n13398_not
g47372 not n19743 ; n19743_not
g47373 not n24396 ; n24396_not
g47374 not n13569 ; n13569_not
g47375 not n24288 ; n24288_not
g47376 not n24468 ; n24468_not
g47377 not n13776 ; n13776_not
g47378 not n24297 ; n24297_not
g47379 not n19905 ; n19905_not
g47380 not n13767 ; n13767_not
g47381 not n23928 ; n23928_not
g47382 not n13947 ; n13947_not
g47383 not n24387 ; n24387_not
g47384 not n10896 ; n10896_not
g47385 not n26367 ; n26367_not
g47386 not n18960 ; n18960_not
g47387 not n26358 ; n26358_not
g47388 not n26286 ; n26286_not
g47389 not n26349 ; n26349_not
g47390 not n18663 ; n18663_not
g47391 not n10959 ; n10959_not
g47392 not n10968 ; n10968_not
g47393 not n10977 ; n10977_not
g47394 not n26187 ; n26187_not
g47395 not n26295 ; n26295_not
g47396 not n10986 ; n10986_not
g47397 not n26277 ; n26277_not
g47398 not n10995 ; n10995_not
g47399 not n26259 ; n26259_not
g47400 not n18690 ; n18690_not
g47401 not n10878 ; n10878_not
g47402 not n18645 ; n18645_not
g47403 not n18636 ; n18636_not
g47404 not n19059 ; n19059_not
g47405 not n26529 ; n26529_not
g47406 not n10788 ; n10788_not
g47407 not n10797 ; n10797_not
g47408 not n26439 ; n26439_not
g47409 not n18915 ; n18915_not
g47410 not n26493 ; n26493_not
g47411 not n26484 ; n26484_not
g47412 not n18924 ; n18924_not
g47413 not n26475 ; n26475_not
g47414 not n10779 ; n10779_not
g47415 not n26457 ; n26457_not
g47416 not n26394 ; n26394_not
g47417 not n26448 ; n26448_not
g47418 not n18942 ; n18942_not
g47419 not n10869 ; n10869_not
g47420 not n18951 ; n18951_not
g47421 not n10887 ; n10887_not
g47422 not n26385 ; n26385_not
g47423 not n25944 ; n25944_not
g47424 not n19158 ; n19158_not
g47425 not n11769 ; n11769_not
g47426 not n11778 ; n11778_not
g47427 not n19167 ; n19167_not
g47428 not n11787 ; n11787_not
g47429 not n11796 ; n11796_not
g47430 not n25755 ; n25755_not
g47431 not n19185 ; n19185_not
g47432 not n11688 ; n11688_not
g47433 not n25935 ; n25935_not
g47434 not n25980 ; n25980_not
g47435 not n25962 ; n25962_not
g47436 not n25953 ; n25953_not
g47437 not n11859 ; n11859_not
g47438 not n25827 ; n25827_not
g47439 not n25926 ; n25926_not
g47440 not n25908 ; n25908_not
g47441 not n19194 ; n19194_not
g47442 not n25854 ; n25854_not
g47443 not n18564 ; n18564_not
g47444 not n25890 ; n25890_not
g47445 not n18861 ; n18861_not
g47446 not n19068 ; n19068_not
g47447 not n18627 ; n18627_not
g47448 not n26196 ; n26196_not
g47449 not n19077 ; n19077_not
g47450 not n26178 ; n26178_not
g47451 not n11499 ; n11499_not
g47452 not n26097 ; n26097_not
g47453 not n19095 ; n19095_not
g47454 not n18780 ; n18780_not
g47455 not n18618 ; n18618_not
g47456 not n11589 ; n11589_not
g47457 not n18609 ; n18609_not
g47458 not n11598 ; n11598_not
g47459 not n18591 ; n18591_not
g47460 not n11679 ; n11679_not
g47461 not n18285 ; n18285_not
g47462 not n19149 ; n19149_not
g47463 not n18582 ; n18582_not
g47464 not n27069 ; n27069_not
g47465 not n26970 ; n26970_not
g47466 not n18492 ; n18492_not
g47467 not n18771 ; n18771_not
g47468 not n26961 ; n26961_not
g47469 not n26952 ; n26952_not
g47470 not n26943 ; n26943_not
g47471 not n26934 ; n26934_not
g47472 not n26925 ; n26925_not
g47473 not n26916 ; n26916_not
g47474 not n18672 ; n18672_not
g47475 not n26907 ; n26907_not
g47476 not n18807 ; n18807_not
g47477 not n26880 ; n26880_not
g47478 not n26871 ; n26871_not
g47479 not n26862 ; n26862_not
g47480 not n26781 ; n26781_not
g47481 not n26853 ; n26853_not
g47482 not n27294 ; n27294_not
g47483 not n27285 ; n27285_not
g47484 not n27267 ; n27267_not
g47485 not n27276 ; n27276_not
g47486 not n18348 ; n18348_not
g47487 not n18708 ; n18708_not
g47488 not n27195 ; n27195_not
g47489 not n18717 ; n18717_not
g47490 not n27186 ; n27186_not
g47491 not n27177 ; n27177_not
g47492 not n27168 ; n27168_not
g47493 not n27159 ; n27159_not
g47494 not n18735 ; n18735_not
g47495 not n27096 ; n27096_not
g47496 not n18744 ; n18744_not
g47497 not n27078 ; n27078_not
g47498 not n27087 ; n27087_not
g47499 not n26619 ; n26619_not
g47500 not n26709 ; n26709_not
g47501 not n18852 ; n18852_not
g47502 not n26637 ; n26637_not
g47503 not n26691 ; n26691_not
g47504 not n26574 ; n26574_not
g47505 not n26565 ; n26565_not
g47506 not n26664 ; n26664_not
g47507 not n26655 ; n26655_not
g47508 not n26592 ; n26592_not
g47509 not n10689 ; n10689_not
g47510 not n26628 ; n26628_not
g47511 not n18870 ; n18870_not
g47512 not n10698 ; n10698_not
g47513 not n26583 ; n26583_not
g47514 not n26556 ; n26556_not
g47515 not n26547 ; n26547_not
g47516 not n26538 ; n26538_not
g47517 not n18906 ; n18906_not
g47518 not n26844 ; n26844_not
g47519 not n26835 ; n26835_not
g47520 not n26826 ; n26826_not
g47521 not n26817 ; n26817_not
g47522 not n18816 ; n18816_not
g47523 not n18825 ; n18825_not
g47524 not n26808 ; n26808_not
g47525 not n26790 ; n26790_not
g47526 not n26772 ; n26772_not
g47527 not n26763 ; n26763_not
g47528 not n26727 ; n26727_not
g47529 not n26754 ; n26754_not
g47530 not n18834 ; n18834_not
g47531 not n26682 ; n26682_not
g47532 not n26736 ; n26736_not
g47533 not n18762 ; n18762_not
g47534 not n10599 ; n10599_not
g47535 not n18843 ; n18843_not
g47536 not n19626 ; n19626_not
g47537 not n12975 ; n12975_not
g47538 not n24981 ; n24981_not
g47539 not n24963 ; n24963_not
g47540 not n24954 ; n24954_not
g47541 not n24783 ; n24783_not
g47542 not n18456 ; n18456_not
g47543 not n24945 ; n24945_not
g47544 not n24936 ; n24936_not
g47545 not n19635 ; n19635_not
g47546 not n24927 ; n24927_not
g47547 not n24918 ; n24918_not
g47548 not n24909 ; n24909_not
g47549 not n19644 ; n19644_not
g47550 not n12984 ; n12984_not
g47551 not n24891 ; n24891_not
g47552 not n24882 ; n24882_not
g47553 not n24873 ; n24873_not
g47554 not n24864 ; n24864_not
g47555 not n24639 ; n24639_not
g47556 not n24855 ; n24855_not
g47557 not n25179 ; n25179_not
g47558 not n19428 ; n19428_not
g47559 not n12768 ; n12768_not
g47560 not n19563 ; n19563_not
g47561 not n12777 ; n12777_not
g47562 not n12786 ; n12786_not
g47563 not n19572 ; n19572_not
g47564 not n25098 ; n25098_not
g47565 not n19590 ; n19590_not
g47566 not n12858 ; n12858_not
g47567 not n25089 ; n25089_not
g47568 not n12867 ; n12867_not
g47569 not n12876 ; n12876_not
g47570 not n24972 ; n24972_not
g47571 not n12885 ; n12885_not
g47572 not n12894 ; n12894_not
g47573 not n19608 ; n19608_not
g47574 not n18465 ; n18465_not
g47575 not n12939 ; n12939_not
g47576 not n19617 ; n19617_not
g47577 not n12966 ; n12966_not
g47578 not n24675 ; n24675_not
g47579 not n24666 ; n24666_not
g47580 not n24657 ; n24657_not
g47581 not n19734 ; n19734_not
g47582 not n24648 ; n24648_not
g47583 not n19752 ; n19752_not
g47584 not n13299 ; n13299_not
g47585 not n24594 ; n24594_not
g47586 not n19770 ; n19770_not
g47587 not n24585 ; n24585_not
g47588 not n13389 ; n13389_not
g47589 not n24567 ; n24567_not
g47590 not n24549 ; n24549_not
g47591 not n19815 ; n19815_not
g47592 not n19527 ; n19527_not
g47593 not n24495 ; n24495_not
g47594 not n24486 ; n24486_not
g47595 not n12993 ; n12993_not
g47596 not n24846 ; n24846_not
g47597 not n19653 ; n19653_not
g47598 not n24828 ; n24828_not
g47599 not n24819 ; n24819_not
g47600 not n24729 ; n24729_not
g47601 not n24792 ; n24792_not
g47602 not n12678 ; n12678_not
g47603 not n24774 ; n24774_not
g47604 not n19671 ; n19671_not
g47605 not n24765 ; n24765_not
g47606 not n24756 ; n24756_not
g47607 not n19680 ; n19680_not
g47608 not n24747 ; n24747_not
g47609 not n24738 ; n24738_not
g47610 not n19707 ; n19707_not
g47611 not n18447 ; n18447_not
g47612 not n19716 ; n19716_not
g47613 not n24693 ; n24693_not
g47614 not n24684 ; n24684_not
g47615 not n19248 ; n19248_not
g47616 not n25728 ; n25728_not
g47617 not n19257 ; n19257_not
g47618 not n18555 ; n18555_not
g47619 not n25719 ; n25719_not
g47620 not n11949 ; n11949_not
g47621 not n25683 ; n25683_not
g47622 not n25674 ; n25674_not
g47623 not n19275 ; n19275_not
g47624 not n19266 ; n19266_not
g47625 not n25665 ; n25665_not
g47626 not n25656 ; n25656_not
g47627 not n25647 ; n25647_not
g47628 not n25638 ; n25638_not
g47629 not n11868 ; n11868_not
g47630 not n25629 ; n25629_not
g47631 not n19293 ; n19293_not
g47632 not n11967 ; n11967_not
g47633 not n11976 ; n11976_not
g47634 not n25593 ; n25593_not
g47635 not n25584 ; n25584_not
g47636 not n25575 ; n25575_not
g47637 not n25881 ; n25881_not
g47638 not n25746 ; n25746_not
g47639 not n25863 ; n25863_not
g47640 not n25872 ; n25872_not
g47641 not n18573 ; n18573_not
g47642 not n25845 ; n25845_not
g47643 not n25782 ; n25782_not
g47644 not n25836 ; n25836_not
g47645 not n11877 ; n11877_not
g47646 not n25818 ; n25818_not
g47647 not n11886 ; n11886_not
g47648 not n25809 ; n25809_not
g47649 not n25791 ; n25791_not
g47650 not n25773 ; n25773_not
g47651 not n25764 ; n25764_not
g47652 not n19239 ; n19239_not
g47653 not n25737 ; n25737_not
g47654 not n19419 ; n19419_not
g47655 not n25395 ; n25395_not
g47656 not n25386 ; n25386_not
g47657 not n25368 ; n25368_not
g47658 not n25377 ; n25377_not
g47659 not n19437 ; n19437_not
g47660 not n12498 ; n12498_not
g47661 not n19455 ; n19455_not
g47662 not n19473 ; n19473_not
g47663 not n12588 ; n12588_not
g47664 not n25296 ; n25296_not
g47665 not n25287 ; n25287_not
g47666 not n12597 ; n12597_not
g47667 not n19491 ; n19491_not
g47668 not n19509 ; n19509_not
g47669 not n18483 ; n18483_not
g47670 not n12669 ; n12669_not
g47671 not n12687 ; n12687_not
g47672 not n12696 ; n12696_not
g47673 not n19536 ; n19536_not
g47674 not n25197 ; n25197_not
g47675 not n25188 ; n25188_not
g47676 not n12759 ; n12759_not
g47677 not n11985 ; n11985_not
g47678 not n25557 ; n25557_not
g47679 not n11994 ; n11994_not
g47680 not n25539 ; n25539_not
g47681 not n25476 ; n25476_not
g47682 not n18537 ; n18537_not
g47683 not n19329 ; n19329_not
g47684 not n19338 ; n19338_not
g47685 not n18528 ; n18528_not
g47686 not n25494 ; n25494_not
g47687 not n19356 ; n19356_not
g47688 not n25485 ; n25485_not
g47689 not n19365 ; n19365_not
g47690 not n25458 ; n25458_not
g47691 not n25449 ; n25449_not
g47692 not n19374 ; n19374_not
g47693 not n19383 ; n19383_not
g47694 not n18519 ; n18519_not
g47695 not n12399 ; n12399_not
g47696 not n22785 ; n22785_not
g47697 not n14937 ; n14937_not
g47698 not n17808 ; n17808_not
g47699 not n22992 ; n22992_not
g47700 not n14982 ; n14982_not
g47701 not n15369 ; n15369_not
g47702 not n22983 ; n22983_not
g47703 not n22974 ; n22974_not
g47704 not n17790 ; n17790_not
g47705 not n22965 ; n22965_not
g47706 not n17781 ; n17781_not
g47707 not n22956 ; n22956_not
g47708 not n22938 ; n22938_not
g47709 not n22893 ; n22893_not
g47710 not n15387 ; n15387_not
g47711 not n22929 ; n22929_not
g47712 not n15396 ; n15396_not
g47713 not n17763 ; n17763_not
g47714 not n14586 ; n14586_not
g47715 not n14991 ; n14991_not
g47716 not n14694 ; n14694_not
g47717 not n17880 ; n17880_not
g47718 not n17871 ; n17871_not
g47719 not n15099 ; n15099_not
g47720 not n14766 ; n14766_not
g47721 not n17862 ; n17862_not
g47722 not n15189 ; n15189_not
g47723 not n17844 ; n17844_not
g47724 not n20499 ; n20499_not
g47725 not n15198 ; n15198_not
g47726 not n14856 ; n14856_not
g47727 not n17835 ; n17835_not
g47728 not n17772 ; n17772_not
g47729 not n17826 ; n17826_not
g47730 not n15279 ; n15279_not
g47731 not n15288 ; n15288_not
g47732 not n17817 ; n17817_not
g47733 not n15297 ; n15297_not
g47734 not n15549 ; n15549_not
g47735 not n15558 ; n15558_not
g47736 not n17673 ; n17673_not
g47737 not n20679 ; n20679_not
g47738 not n15567 ; n15567_not
g47739 not n15576 ; n15576_not
g47740 not n22695 ; n22695_not
g47741 not n17664 ; n17664_not
g47742 not n22686 ; n22686_not
g47743 not n22677 ; n22677_not
g47744 not n15585 ; n15585_not
g47745 not n22668 ; n22668_not
g47746 not n20697 ; n20697_not
g47747 not n22659 ; n22659_not
g47748 not n17655 ; n17655_not
g47749 not n17646 ; n17646_not
g47750 not n17637 ; n17637_not
g47751 not n17628 ; n17628_not
g47752 not n15648 ; n15648_not
g47753 not n15666 ; n15666_not
g47754 not n15495 ; n15495_not
g47755 not n22596 ; n22596_not
g47756 not n22875 ; n22875_not
g47757 not n22884 ; n22884_not
g47758 not n22866 ; n22866_not
g47759 not n17754 ; n17754_not
g47760 not n22848 ; n22848_not
g47761 not n22839 ; n22839_not
g47762 not n20598 ; n20598_not
g47763 not n15468 ; n15468_not
g47764 not n15477 ; n15477_not
g47765 not n17457 ; n17457_not
g47766 not n17745 ; n17745_not
g47767 not n15486 ; n15486_not
g47768 not n17727 ; n17727_not
g47769 not n17718 ; n17718_not
g47770 not n17529 ; n17529_not
g47771 not n22794 ; n22794_not
g47772 not n22479 ; n22479_not
g47773 not n17691 ; n17691_not
g47774 not n22758 ; n22758_not
g47775 not n22767 ; n22767_not
g47776 not n22488 ; n22488_not
g47777 not n22749 ; n22749_not
g47778 not n17682 ; n17682_not
g47779 not n14595 ; n14595_not
g47780 not n23577 ; n23577_not
g47781 not n23586 ; n23586_not
g47782 not n19941 ; n19941_not
g47783 not n23568 ; n23568_not
g47784 not n18096 ; n18096_not
g47785 not n23559 ; n23559_not
g47786 not n23397 ; n23397_not
g47787 not n18078 ; n18078_not
g47788 not n14649 ; n14649_not
g47789 not n14658 ; n14658_not
g47790 not n14667 ; n14667_not
g47791 not n17907 ; n17907_not
g47792 not n14676 ; n14676_not
g47793 not n14685 ; n14685_not
g47794 not n23496 ; n23496_not
g47795 not n18267 ; n18267_not
g47796 not n17916 ; n17916_not
g47797 not n18258 ; n18258_not
g47798 not n14496 ; n14496_not
g47799 not n18249 ; n18249_not
g47800 not n23658 ; n23658_not
g47801 not n23685 ; n23685_not
g47802 not n23694 ; n23694_not
g47803 not n23676 ; n23676_not
g47804 not n23667 ; n23667_not
g47805 not n18195 ; n18195_not
g47806 not n18186 ; n18186_not
g47807 not n23649 ; n23649_not
g47808 not n23469 ; n23469_not
g47809 not n14559 ; n14559_not
g47810 not n18177 ; n18177_not
g47811 not n18168 ; n18168_not
g47812 not n14577 ; n14577_not
g47813 not n14568 ; n14568_not
g47814 not n18159 ; n18159_not
g47815 not n17943 ; n17943_not
g47816 not n14865 ; n14865_not
g47817 not n14874 ; n14874_not
g47818 not n14883 ; n14883_not
g47819 not n23298 ; n23298_not
g47820 not n17934 ; n17934_not
g47821 not n14892 ; n14892_not
g47822 not n17709 ; n17709_not
g47823 not n14928 ; n14928_not
g47824 not n17736 ; n17736_not
g47825 not n14946 ; n14946_not
g47826 not n14955 ; n14955_not
g47827 not n14964 ; n14964_not
g47828 not n23199 ; n23199_not
g47829 not n14973 ; n14973_not
g47830 not n23487 ; n23487_not
g47831 not n23478 ; n23478_not
g47832 not n17952 ; n17952_not
g47833 not n14739 ; n14739_not
g47834 not n14748 ; n14748_not
g47835 not n14757 ; n14757_not
g47836 not n14775 ; n14775_not
g47837 not n14784 ; n14784_not
g47838 not n14298 ; n14298_not
g47839 not n23388 ; n23388_not
g47840 not n14793 ; n14793_not
g47841 not n23379 ; n23379_not
g47842 not n17961 ; n17961_not
g47843 not n14829 ; n14829_not
g47844 not n14838 ; n14838_not
g47845 not n14847 ; n14847_not
g47846 not n16575 ; n16575_not
g47847 not n21786 ; n21786_not
g47848 not n21777 ; n21777_not
g47849 not n16584 ; n16584_not
g47850 not n21768 ; n21768_not
g47851 not n17268 ; n17268_not
g47852 not n16467 ; n16467_not
g47853 not n21759 ; n21759_not
g47854 not n20859 ; n20859_not
g47855 not n17259 ; n17259_not
g47856 not n16368 ; n16368_not
g47857 not n21489 ; n21489_not
g47858 not n16908 ; n16908_not
g47859 not n16638 ; n16638_not
g47860 not n16647 ; n16647_not
g47861 not n16656 ; n16656_not
g47862 not n16665 ; n16665_not
g47863 not n21678 ; n21678_not
g47864 not n21687 ; n21687_not
g47865 not n16629 ; n16629_not
g47866 not n16674 ; n16674_not
g47867 not n21975 ; n21975_not
g47868 not n21966 ; n21966_not
g47869 not n16458 ; n16458_not
g47870 not n17394 ; n17394_not
g47871 not n21939 ; n21939_not
g47872 not n16476 ; n16476_not
g47873 not n16485 ; n16485_not
g47874 not n17367 ; n17367_not
g47875 not n21894 ; n21894_not
g47876 not n21876 ; n21876_not
g47877 not n21867 ; n21867_not
g47878 not n21858 ; n21858_not
g47879 not n17349 ; n17349_not
g47880 not n16539 ; n16539_not
g47881 not n16548 ; n16548_not
g47882 not n16557 ; n16557_not
g47883 not n17295 ; n17295_not
g47884 not n17286 ; n17286_not
g47885 not n16818 ; n16818_not
g47886 not n16827 ; n16827_not
g47887 not n21498 ; n21498_not
g47888 not n16836 ; n16836_not
g47889 not n16854 ; n16854_not
g47890 not n16863 ; n16863_not
g47891 not n16872 ; n16872_not
g47892 not n16881 ; n16881_not
g47893 not n21399 ; n21399_not
g47894 not n16917 ; n16917_not
g47895 not n16971 ; n16971_not
g47896 not n16926 ; n16926_not
g47897 not n16980 ; n16980_not
g47898 not n16935 ; n16935_not
g47899 not n16953 ; n16953_not
g47900 not n16962 ; n16962_not
g47901 not n16809 ; n16809_not
g47902 not n21669 ; n21669_not
g47903 not n16683 ; n16683_not
g47904 not n17196 ; n17196_not
g47905 not n16692 ; n16692_not
g47906 not n17187 ; n17187_not
g47907 not n16719 ; n16719_not
g47908 not n17178 ; n17178_not
g47909 not n16737 ; n16737_not
g47910 not n16746 ; n16746_not
g47911 not n16755 ; n16755_not
g47912 not n21597 ; n21597_not
g47913 not n21588 ; n21588_not
g47914 not n16764 ; n16764_not
g47915 not n21579 ; n21579_not
g47916 not n17097 ; n17097_not
g47917 not n17088 ; n17088_not
g47918 not n16782 ; n16782_not
g47919 not n16791 ; n16791_not
g47920 not n17079 ; n17079_not
g47921 not n17565 ; n17565_not
g47922 not n15828 ; n15828_not
g47923 not n15846 ; n15846_not
g47924 not n17556 ; n17556_not
g47925 not n22398 ; n22398_not
g47926 not n22389 ; n22389_not
g47927 not n15855 ; n15855_not
g47928 not n15882 ; n15882_not
g47929 not n15891 ; n15891_not
g47930 not n17547 ; n17547_not
g47931 not n15909 ; n15909_not
g47932 not n17538 ; n17538_not
g47933 not n15927 ; n15927_not
g47934 not n20868 ; n20868_not
g47935 not n15936 ; n15936_not
g47936 not n22299 ; n22299_not
g47937 not n15945 ; n15945_not
g47938 not n22587 ; n22587_not
g47939 not n22578 ; n22578_not
g47940 not n17592 ; n17592_not
g47941 not n15684 ; n15684_not
g47942 not n22569 ; n22569_not
g47943 not n15675 ; n15675_not
g47944 not n15693 ; n15693_not
g47945 not n20769 ; n20769_not
g47946 not n20778 ; n20778_not
g47947 not n15729 ; n15729_not
g47948 not n15738 ; n15738_not
g47949 not n15747 ; n15747_not
g47950 not n15756 ; n15756_not
g47951 not n15378 ; n15378_not
g47952 not n20796 ; n20796_not
g47953 not n20787 ; n20787_not
g47954 not n17583 ; n17583_not
g47955 not n15783 ; n15783_not
g47956 not n15792 ; n15792_not
g47957 not n15819 ; n15819_not
g47958 not n16269 ; n16269_not
g47959 not n20967 ; n20967_not
g47960 not n16278 ; n16278_not
g47961 not n16287 ; n16287_not
g47962 not n15864 ; n15864_not
g47963 not n16296 ; n16296_not
g47964 not n20985 ; n20985_not
g47965 not n20976 ; n20976_not
g47966 not n16359 ; n16359_not
g47967 not n20994 ; n20994_not
g47968 not n17466 ; n17466_not
g47969 not n16377 ; n16377_not
g47970 not n16386 ; n16386_not
g47971 not n16395 ; n16395_not
g47972 not n17448 ; n17448_not
g47973 not n16449 ; n16449_not
g47974 not n21993 ; n21993_not
g47975 not n21984 ; n21984_not
g47976 not n15954 ; n15954_not
g47977 not n20886 ; n20886_not
g47978 not n15963 ; n15963_not
g47979 not n15972 ; n15972_not
g47980 not n15981 ; n15981_not
g47981 not n15990 ; n15990_not
g47982 not n21885 ; n21885_not
g47983 not n20895 ; n20895_not
g47984 not n17358 ; n17358_not
g47985 not n16089 ; n16089_not
g47986 not n16098 ; n16098_not
g47987 not n17493 ; n17493_not
g47988 not n17484 ; n17484_not
g47989 not n21957 ; n21957_not
g47990 not n16197 ; n16197_not
g47991 not n20949 ; n20949_not
g47992 not n17475 ; n17475_not
g47993 not n20958 ; n20958_not
g47994 not n18375 ; n18375_not
g47995 not n23892 ; n23892_not
g47996 not n14379 ; n14379_not
g47997 not n23748 ; n23748_not
g47998 not n18276 ; n18276_not
g47999 not n14388 ; n14388_not
g48000 not n23775 ; n23775_not
g48001 not n23937 ; n23937_not
g48002 not n14397 ; n14397_not
g48003 not n23766 ; n23766_not
g48004 not n14478 ; n14478_not
g48005 not n18294 ; n18294_not
g48006 not n23874 ; n23874_not
g48007 not n23964 ; n23964_not
g48008 not n23793 ; n23793_not
g48009 not n23865 ; n23865_not
g48010 not n23955 ; n23955_not
g48011 not n23757 ; n23757_not
g48012 not n23784 ; n23784_not
g48013 not n23838 ; n23838_not
g48014 not n14469 ; n14469_not
g48015 not n23847 ; n23847_not
g48016 not n23982 ; n23982_not
g48017 not n23919 ; n23919_not
g48018 not n23595 ; n23595_not
g48019 not n23739 ; n23739_not
g48020 not n14289 ; n14289_not
g48021 not n18357 ; n18357_not
g48022 not n18393 ; n18393_not
g48023 not n18366 ; n18366_not
g48024 not n19285 ; n19285_not
g48025 not n17287 ; n17287_not
g48026 not n25639 ; n25639_not
g48027 not n19069 ; n19069_not
g48028 not n11959 ; n11959_not
g48029 not n25495 ; n25495_not
g48030 not n15595 ; n15595_not
g48031 not n25558 ; n25558_not
g48032 not n20698 ; n20698_not
g48033 not n13876 ; n13876_not
g48034 not n23884 ; n23884_not
g48035 not n22669 ; n22669_not
g48036 not n15586 ; n15586_not
g48037 not n15667 ; n15667_not
g48038 not n25675 ; n25675_not
g48039 not n15649 ; n15649_not
g48040 not n19276 ; n19276_not
g48041 not n19195 ; n19195_not
g48042 not n25666 ; n25666_not
g48043 not n17629 ; n17629_not
g48044 not n18358 ; n18358_not
g48045 not n17548 ; n17548_not
g48046 not n13885 ; n13885_not
g48047 not n19933 ; n19933_not
g48048 not n25657 ; n25657_not
g48049 not n17647 ; n17647_not
g48050 not n25648 ; n25648_not
g48051 not n17656 ; n17656_not
g48052 not n25585 ; n25585_not
g48053 not n25576 ; n25576_not
g48054 not n15577 ; n15577_not
g48055 not n18673 ; n18673_not
g48056 not n25567 ; n25567_not
g48057 not n25972 ; n25972_not
g48058 not n25936 ; n25936_not
g48059 not n11986 ; n11986_not
g48060 not n15568 ; n15568_not
g48061 not n13867 ; n13867_not
g48062 not n23866 ; n23866_not
g48063 not n17674 ; n17674_not
g48064 not n18547 ; n18547_not
g48065 not n15559 ; n15559_not
g48066 not n11968 ; n11968_not
g48067 not n22678 ; n22678_not
g48068 not n17665 ; n17665_not
g48069 not n19294 ; n19294_not
g48070 not n15874 ; n15874_not
g48071 not n25945 ; n25945_not
g48072 not n22687 ; n22687_not
g48073 not n25954 ; n25954_not
g48074 not n11977 ; n11977_not
g48075 not n20689 ; n20689_not
g48076 not n25594 ; n25594_not
g48077 not n25963 ; n25963_not
g48078 not n22696 ; n22696_not
g48079 not n15766 ; n15766_not
g48080 not n25819 ; n25819_not
g48081 not n17584 ; n17584_not
g48082 not n25882 ; n25882_not
g48083 not n11878 ; n11878_not
g48084 not n25891 ; n25891_not
g48085 not n18565 ; n18565_not
g48086 not n20797 ; n20797_not
g48087 not n11887 ; n11887_not
g48088 not n17557 ; n17557_not
g48089 not n22399 ; n22399_not
g48090 not n25792 ; n25792_not
g48091 not n22489 ; n22489_not
g48092 not n15757 ; n15757_not
g48093 not n25783 ; n25783_not
g48094 not n20788 ; n20788_not
g48095 not n18349 ; n18349_not
g48096 not n17575 ; n17575_not
g48097 not n25864 ; n25864_not
g48098 not n11869 ; n11869_not
g48099 not n25855 ; n25855_not
g48100 not n18574 ; n18574_not
g48101 not n15793 ; n15793_not
g48102 not n25873 ; n25873_not
g48103 not n25846 ; n25846_not
g48104 not n15784 ; n15784_not
g48105 not n25837 ; n25837_not
g48106 not n25828 ; n25828_not
g48107 not n15829 ; n15829_not
g48108 not n15838 ; n15838_not
g48109 not n17593 ; n17593_not
g48110 not n15694 ; n15694_not
g48111 not n25729 ; n25729_not
g48112 not n19258 ; n19258_not
g48113 not n15676 ; n15676_not
g48114 not n15685 ; n15685_not
g48115 not n23893 ; n23893_not
g48116 not n22579 ; n22579_not
g48117 not n18925 ; n18925_not
g48118 not n25927 ; n25927_not
g48119 not n19267 ; n19267_not
g48120 not n25693 ; n25693_not
g48121 not n22597 ; n22597_not
g48122 not n24199 ; n24199_not
g48123 not n25684 ; n25684_not
g48124 not n15748 ; n15748_not
g48125 not n25765 ; n25765_not
g48126 not n25756 ; n25756_not
g48127 not n25909 ; n25909_not
g48128 not n15739 ; n15739_not
g48129 not n25747 ; n25747_not
g48130 not n25918 ; n25918_not
g48131 not n20779 ; n20779_not
g48132 not n15856 ; n15856_not
g48133 not n18556 ; n18556_not
g48134 not n25738 ; n25738_not
g48135 not n19249 ; n19249_not
g48136 not n12688 ; n12688_not
g48137 not n14389 ; n14389_not
g48138 not n12697 ; n12697_not
g48139 not n17836 ; n17836_not
g48140 not n19537 ; n19537_not
g48141 not n19546 ; n19546_not
g48142 not n25198 ; n25198_not
g48143 not n15199 ; n15199_not
g48144 not n14398 ; n14398_not
g48145 not n25189 ; n25189_not
g48146 not n17845 ; n17845_not
g48147 not n22966 ; n22966_not
g48148 not n19555 ; n19555_not
g48149 not n14785 ; n14785_not
g48150 not n17863 ; n17863_not
g48151 not n17476 ; n17476_not
g48152 not n12769 ; n12769_not
g48153 not n17971 ; n17971_not
g48154 not n22993 ; n22993_not
g48155 not n12589 ; n12589_not
g48156 not n25279 ; n25279_not
g48157 not n25288 ; n25288_not
g48158 not n12598 ; n12598_not
g48159 not n19492 ; n19492_not
g48160 not n14965 ; n14965_not
g48161 not n17809 ; n17809_not
g48162 not n18484 ; n18484_not
g48163 not n15298 ; n15298_not
g48164 not n15289 ; n15289_not
g48165 not n13786 ; n13786_not
g48166 not n12679 ; n12679_not
g48167 not n17827 ; n17827_not
g48168 not n19528 ; n19528_not
g48169 not n18475 ; n18475_not
g48170 not n17818 ; n17818_not
g48171 not n12895 ; n12895_not
g48172 not n14974 ; n14974_not
g48173 not n24865 ; n24865_not
g48174 not n19609 ; n19609_not
g48175 not n18466 ; n18466_not
g48176 not n24289 ; n24289_not
g48177 not n12949 ; n12949_not
g48178 not n17890 ; n17890_not
g48179 not n12958 ; n12958_not
g48180 not n14956 ; n14956_not
g48181 not n12967 ; n12967_not
g48182 not n13777 ; n13777_not
g48183 not n19627 ; n19627_not
g48184 not n14947 ; n14947_not
g48185 not n24982 ; n24982_not
g48186 not n12976 ; n12976_not
g48187 not n19564 ; n19564_not
g48188 not n12778 ; n12778_not
g48189 not n14749 ; n14749_not
g48190 not n12787 ; n12787_not
g48191 not n12796 ; n12796_not
g48192 not n24793 ; n24793_not
g48193 not n17881 ; n17881_not
g48194 not n19582 ; n19582_not
g48195 not n25099 ; n25099_not
g48196 not n24928 ; n24928_not
g48197 not n19591 ; n19591_not
g48198 not n14992 ; n14992_not
g48199 not n12859 ; n12859_not
g48200 not n14983 ; n14983_not
g48201 not n12877 ; n12877_not
g48202 not n24973 ; n24973_not
g48203 not n12886 ; n12886_not
g48204 not n17719 ; n17719_not
g48205 not n25477 ; n25477_not
g48206 not n15487 ; n15487_not
g48207 not n17737 ; n17737_not
g48208 not n15478 ; n15478_not
g48209 not n17746 ; n17746_not
g48210 not n19366 ; n19366_not
g48211 not n25459 ; n25459_not
g48212 not n20599 ; n20599_not
g48213 not n23848 ; n23848_not
g48214 not n22849 ; n22849_not
g48215 not n17755 ; n17755_not
g48216 not n19375 ; n19375_not
g48217 not n23668 ; n23668_not
g48218 not n22858 ; n22858_not
g48219 not n25549 ; n25549_not
g48220 not n11995 ; n11995_not
g48221 not n13858 ; n13858_not
g48222 not n17683 ; n17683_not
g48223 not n13678 ; n13678_not
g48224 not n22759 ; n22759_not
g48225 not n23875 ; n23875_not
g48226 not n18538 ; n18538_not
g48227 not n22768 ; n22768_not
g48228 not n22777 ; n22777_not
g48229 not n17692 ; n17692_not
g48230 not n19339 ; n19339_not
g48231 not n22786 ; n22786_not
g48232 not n18439 ; n18439_not
g48233 not n22795 ; n22795_not
g48234 not n18529 ; n18529_not
g48235 not n15496 ; n15496_not
g48236 not n25486 ; n25486_not
g48237 not n22939 ; n22939_not
g48238 not n15379 ; n15379_not
g48239 not n17773 ; n17773_not
g48240 not n19447 ; n19447_not
g48241 not n22957 ; n22957_not
g48242 not n17782 ; n17782_not
g48243 not n19078 ; n19078_not
g48244 not n19456 ; n19456_not
g48245 not n12499 ; n12499_not
g48246 not n22975 ; n22975_not
g48247 not n17791 ; n17791_not
g48248 not n19474 ; n19474_not
g48249 not n22984 ; n22984_not
g48250 not n19483 ; n19483_not
g48251 not n25297 ; n25297_not
g48252 not n22867 ; n22867_not
g48253 not n22876 ; n22876_not
g48254 not n19384 ; n19384_not
g48255 not n22885 ; n22885_not
g48256 not n22894 ; n22894_not
g48257 not n25396 ; n25396_not
g48258 not n15397 ; n15397_not
g48259 not n25387 ; n25387_not
g48260 not n19429 ; n19429_not
g48261 not n19924 ; n19924_not
g48262 not n25378 ; n25378_not
g48263 not n15388 ; n15388_not
g48264 not n23839 ; n23839_not
g48265 not n25369 ; n25369_not
g48266 not n19438 ; n19438_not
g48267 not n26746 ; n26746_not
g48268 not n26683 ; n26683_not
g48269 not n18835 ; n18835_not
g48270 not n16684 ; n16684_not
g48271 not n26737 ; n26737_not
g48272 not n17197 ; n17197_not
g48273 not n23974 ; n23974_not
g48274 not n26728 ; n26728_not
g48275 not n16675 ; n16675_not
g48276 not n18844 ; n18844_not
g48277 not n21679 ; n21679_not
g48278 not n21688 ; n21688_not
g48279 not n26629 ; n26629_not
g48280 not n18853 ; n18853_not
g48281 not n16666 ; n16666_not
g48282 not n26692 ; n26692_not
g48283 not n26674 ; n26674_not
g48284 not n16459 ; n16459_not
g48285 not n26818 ; n26818_not
g48286 not n16756 ; n16756_not
g48287 not n18826 ; n18826_not
g48288 not n16738 ; n16738_not
g48289 not n26809 ; n26809_not
g48290 not n17179 ; n17179_not
g48291 not n26791 ; n26791_not
g48292 not n26782 ; n26782_not
g48293 not n17188 ; n17188_not
g48294 not n26773 ; n26773_not
g48295 not n26764 ; n26764_not
g48296 not n23983 ; n23983_not
g48297 not n26755 ; n26755_not
g48298 not n16693 ; n16693_not
g48299 not n26575 ; n26575_not
g48300 not n26476 ; n26476_not
g48301 not n16576 ; n16576_not
g48302 not n26467 ; n26467_not
g48303 not n21769 ; n21769_not
g48304 not n26566 ; n26566_not
g48305 not n26557 ; n26557_not
g48306 not n21796 ; n21796_not
g48307 not n16477 ; n16477_not
g48308 not n26548 ; n26548_not
g48309 not n26539 ; n26539_not
g48310 not n16567 ; n16567_not
g48311 not n17296 ; n17296_not
g48312 not n18907 ; n18907_not
g48313 not n16558 ; n16558_not
g48314 not n16549 ; n16549_not
g48315 not n10789 ; n10789_not
g48316 not n16657 ; n16657_not
g48317 not n21589 ; n21589_not
g48318 not n16648 ; n16648_not
g48319 not n26665 ; n26665_not
g48320 not n26656 ; n26656_not
g48321 not n16891 ; n16891_not
g48322 not n26647 ; n26647_not
g48323 not n20887 ; n20887_not
g48324 not n16387 ; n16387_not
g48325 not n18862 ; n18862_not
g48326 not n16594 ; n16594_not
g48327 not n17269 ; n17269_not
g48328 not n18871 ; n18871_not
g48329 not n10699 ; n10699_not
g48330 not n16585 ; n16585_not
g48331 not n18880 ; n18880_not
g48332 not n26593 ; n26593_not
g48333 not n21778 ; n21778_not
g48334 not n16918 ; n16918_not
g48335 not n13993 ; n13993_not
g48336 not n16909 ; n16909_not
g48337 not n27178 ; n27178_not
g48338 not n16990 ; n16990_not
g48339 not n27097 ; n27097_not
g48340 not n27088 ; n27088_not
g48341 not n16873 ; n16873_not
g48342 not n27079 ; n27079_not
g48343 not n18745 ; n18745_not
g48344 not n18394 ; n18394_not
g48345 not n18754 ; n18754_not
g48346 not n16495 ; n16495_not
g48347 not n18682 ; n18682_not
g48348 not n18763 ; n18763_not
g48349 not n16855 ; n16855_not
g48350 not n19771 ; n19771_not
g48351 not n18772 ; n18772_not
g48352 not n18448 ; n18448_not
g48353 not n27295 ; n27295_not
g48354 not n16963 ; n16963_not
g48355 not n27286 ; n27286_not
g48356 not n23992 ; n23992_not
g48357 not n27268 ; n27268_not
g48358 not n27277 ; n27277_not
g48359 not n16954 ; n16954_not
g48360 not n27259 ; n27259_not
g48361 not n16972 ; n16972_not
g48362 not n16936 ; n16936_not
g48363 not n18709 ; n18709_not
g48364 not n16837 ; n16837_not
g48365 not n27187 ; n27187_not
g48366 not n16981 ; n16981_not
g48367 not n16927 ; n16927_not
g48368 not n18718 ; n18718_not
g48369 not n26908 ; n26908_not
g48370 not n18808 ; n18808_not
g48371 not n26890 ; n26890_not
g48372 not n16792 ; n16792_not
g48373 not n26881 ; n26881_not
g48374 not n23776 ; n23776_not
g48375 not n26872 ; n26872_not
g48376 not n18169 ; n18169_not
g48377 not n26854 ; n26854_not
g48378 not n17089 ; n17089_not
g48379 not n26845 ; n26845_not
g48380 not n26836 ; n26836_not
g48381 not n16765 ; n16765_not
g48382 not n17098 ; n17098_not
g48383 not n18817 ; n18817_not
g48384 not n18781 ; n18781_not
g48385 not n18790 ; n18790_not
g48386 not n26980 ; n26980_not
g48387 not n26971 ; n26971_not
g48388 not n16846 ; n16846_not
g48389 not n26962 ; n26962_not
g48390 not n26935 ; n26935_not
g48391 not n26944 ; n26944_not
g48392 not n26953 ; n26953_not
g48393 not n16639 ; n16639_not
g48394 not n21499 ; n21499_not
g48395 not n16828 ; n16828_not
g48396 not n26926 ; n26926_not
g48397 not n16819 ; n16819_not
g48398 not n26188 ; n26188_not
g48399 not n16198 ; n16198_not
g48400 not n16189 ; n16189_not
g48401 not n17485 ; n17485_not
g48402 not n26179 ; n26179_not
g48403 not n19087 ; n19087_not
g48404 not n26089 ; n26089_not
g48405 not n13957 ; n13957_not
g48406 not n17494 ; n17494_not
g48407 not n16099 ; n16099_not
g48408 not n19096 ; n19096_not
g48409 not n18619 ; n18619_not
g48410 not n13948 ; n13948_not
g48411 not n15847 ; n15847_not
g48412 not n20896 ; n20896_not
g48413 not n15865 ; n15865_not
g48414 not n18637 ; n18637_not
g48415 not n18646 ; n18646_not
g48416 not n20986 ; n20986_not
g48417 not n16297 ; n16297_not
g48418 not n18376 ; n18376_not
g48419 not n20977 ; n20977_not
g48420 not n16288 ; n16288_not
g48421 not n10969 ; n10969_not
g48422 not n16279 ; n16279_not
g48423 not n18628 ; n18628_not
g48424 not n20968 ; n20968_not
g48425 not n23929 ; n23929_not
g48426 not n13966 ; n13966_not
g48427 not n20959 ; n20959_not
g48428 not n26197 ; n26197_not
g48429 not n23938 ; n23938_not
g48430 not n19942 ; n19942_not
g48431 not n17539 ; n17539_not
g48432 not n20869 ; n20869_not
g48433 not n11779 ; n11779_not
g48434 not n19168 ; n19168_not
g48435 not n11788 ; n11788_not
g48436 not n15928 ; n15928_not
g48437 not n19951 ; n19951_not
g48438 not n11797 ; n11797_not
g48439 not n19177 ; n19177_not
g48440 not n15892 ; n15892_not
g48441 not n14299 ; n14299_not
g48442 not n19186 ; n19186_not
g48443 not n25990 ; n25990_not
g48444 not n15883 ; n15883_not
g48445 not n25981 ; n25981_not
g48446 not n11599 ; n11599_not
g48447 not n18592 ; n18592_not
g48448 not n19960 ; n19960_not
g48449 not n26098 ; n26098_not
g48450 not n15982 ; n15982_not
g48451 not n11689 ; n11689_not
g48452 not n18583 ; n18583_not
g48453 not n18367 ; n18367_not
g48454 not n15973 ; n15973_not
g48455 not n15964 ; n15964_not
g48456 not n13939 ; n13939_not
g48457 not n15955 ; n15955_not
g48458 not n19159 ; n19159_not
g48459 not n15946 ; n15946_not
g48460 not n26395 ; n26395_not
g48461 not n26449 ; n26449_not
g48462 not n17368 ; n17368_not
g48463 not n17377 ; n17377_not
g48464 not n16486 ; n16486_not
g48465 not n17386 ; n17386_not
g48466 not n16468 ; n16468_not
g48467 not n10879 ; n10879_not
g48468 not n18952 ; n18952_not
g48469 not n23956 ; n23956_not
g48470 not n17395 ; n17395_not
g48471 not n21949 ; n21949_not
g48472 not n18961 ; n18961_not
g48473 not n26386 ; n26386_not
g48474 not n10798 ; n10798_not
g48475 not n21859 ; n21859_not
g48476 not n18916 ; n18916_not
g48477 not n17359 ; n17359_not
g48478 not n26485 ; n26485_not
g48479 not n21877 ; n21877_not
g48480 not n21868 ; n21868_not
g48481 not n26368 ; n26368_not
g48482 not n21886 ; n21886_not
g48483 not n21895 ; n21895_not
g48484 not n26458 ; n26458_not
g48485 not n10978 ; n10978_not
g48486 not n26296 ; n26296_not
g48487 not n16396 ; n16396_not
g48488 not n13984 ; n13984_not
g48489 not n18655 ; n18655_not
g48490 not n10987 ; n10987_not
g48491 not n26278 ; n26278_not
g48492 not n10996 ; n10996_not
g48493 not n26269 ; n26269_not
g48494 not n16378 ; n16378_not
g48495 not n13975 ; n13975_not
g48496 not n23947 ; n23947_not
g48497 not n17467 ; n17467_not
g48498 not n20995 ; n20995_not
g48499 not n26377 ; n26377_not
g48500 not n10897 ; n10897_not
g48501 not n21958 ; n21958_not
g48502 not n21967 ; n21967_not
g48503 not n18970 ; n18970_not
g48504 not n21976 ; n21976_not
g48505 not n26359 ; n26359_not
g48506 not n26287 ; n26287_not
g48507 not n21985 ; n21985_not
g48508 not n18664 ; n18664_not
g48509 not n17449 ; n17449_not
g48510 not n14569 ; n14569_not
g48511 not n19825 ; n19825_not
g48512 not n24856 ; n24856_not
g48513 not n13687 ; n13687_not
g48514 not n14578 ; n14578_not
g48515 not n24487 ; n24487_not
g48516 not n19744 ; n19744_not
g48517 not n14767 ; n14767_not
g48518 not n24937 ; n24937_not
g48519 not n14587 ; n14587_not
g48520 not n17980 ; n17980_not
g48521 not n23749 ; n23749_not
g48522 not n24748 ; n24748_not
g48523 not n23596 ; n23596_not
g48524 not n18277 ; n18277_not
g48525 not n19816 ; n19816_not
g48526 not n19717 ; n19717_not
g48527 not n24694 ; n24694_not
g48528 not n19807 ; n19807_not
g48529 not n13696 ; n13696_not
g48530 not n14893 ; n14893_not
g48531 not n19843 ; n19843_not
g48532 not n19906 ; n19906_not
g48533 not n24946 ; n24946_not
g48534 not n12994 ; n12994_not
g48535 not n13579 ; n13579_not
g48536 not n23659 ; n23659_not
g48537 not n18196 ; n18196_not
g48538 not n14839 ; n14839_not
g48539 not n17944 ; n17944_not
g48540 not n23794 ; n23794_not
g48541 not n18457 ; n18457_not
g48542 not n24739 ; n24739_not
g48543 not n24298 ; n24298_not
g48544 not n24847 ; n24847_not
g48545 not n18187 ; n18187_not
g48546 not n19834 ; n19834_not
g48547 not n24469 ; n24469_not
g48548 not n19690 ; n19690_not
g48549 not n13768 ; n13768_not
g48550 not n14857 ; n14857_not
g48551 not n18178 ; n18178_not
g48552 not n17926 ; n17926_not
g48553 not n23479 ; n23479_not
g48554 not n14695 ; n14695_not
g48555 not n24568 ; n24568_not
g48556 not n24658 ; n24658_not
g48557 not n14875 ; n14875_not
g48558 not n12985 ; n12985_not
g48559 not n23497 ; n23497_not
g48560 not n23398 ; n23398_not
g48561 not n23758 ; n23758_not
g48562 not n19753 ; n19753_not
g48563 not n18079 ; n18079_not
g48564 not n14479 ; n14479_not
g48565 not n24586 ; n24586_not
g48566 not n24883 ; n24883_not
g48567 not n14677 ; n14677_not
g48568 not n19645 ; n19645_not
g48569 not n14659 ; n14659_not
g48570 not n24595 ; n24595_not
g48571 not n14668 ; n14668_not
g48572 not n24892 ; n24892_not
g48573 not n18286 ; n18286_not
g48574 not n19636 ; n19636_not
g48575 not n13399 ; n13399_not
g48576 not n14866 ; n14866_not
g48577 not n24919 ; n24919_not
g48578 not n24685 ; n24685_not
g48579 not n23587 ; n23587_not
g48580 not n23578 ; n23578_not
g48581 not n24676 ; n24676_not
g48582 not n24874 ; n24874_not
g48583 not n19726 ; n19726_not
g48584 not n17935 ; n17935_not
g48585 not n24667 ; n24667_not
g48586 not n18097 ; n18097_not
g48587 not n19780 ; n19780_not
g48588 not n23767 ; n23767_not
g48589 not n14884 ; n14884_not
g48590 not n19735 ; n19735_not
g48591 not n24559 ; n24559_not
g48592 not n14488 ; n14488_not
g48593 not n24649 ; n24649_not
g48594 not n17917 ; n17917_not
g48595 not n23785 ; n23785_not
g48596 not n19852 ; n19852_not
g48597 not n24784 ; n24784_not
g48598 not n17953 ; n17953_not
g48599 not n19654 ; n19654_not
g48600 not n14497 ; n14497_not
g48601 not n24775 ; n24775_not
g48602 not n18259 ; n18259_not
g48603 not n18268 ; n18268_not
g48604 not n24964 ; n24964_not
g48605 not n19861 ; n19861_not
g48606 not n23695 ; n23695_not
g48607 not n24829 ; n24829_not
g48608 not n13669 ; n13669_not
g48609 not n19672 ; n19672_not
g48610 not n24766 ; n24766_not
g48611 not n13597 ; n13597_not
g48612 not n17962 ; n17962_not
g48613 not n24955 ; n24955_not
g48614 not n14938 ; n14938_not
g48615 not n14794 ; n14794_not
g48616 not n23389 ; n23389_not
g48617 not n19681 ; n19681_not
g48618 not n13588 ; n13588_not
g48619 not n17908 ; n17908_not
g48620 not n24397 ; n24397_not
g48621 not n23677 ; n23677_not
g48622 not n19663 ; n19663_not
g48623 not n23686 ; n23686_not
g48624 not n24379 ; n24379_not
g48625 not n24757 ; n24757_not
g48626 not n15947 ; n15947_not
g48627 not n24785 ; n24785_not
g48628 not n11978 ; n11978_not
g48629 not n18836 ; n18836_not
g48630 not n25595 ; n25595_not
g48631 not n15965 ; n15965_not
g48632 not n17990 ; n17990_not
g48633 not n11699 ; n11699_not
g48634 not n18584 ; n18584_not
g48635 not n19286 ; n19286_not
g48636 not n20699 ; n20699_not
g48637 not n24686 ; n24686_not
g48638 not n23786 ; n23786_not
g48639 not n15893 ; n15893_not
g48640 not n14795 ; n14795_not
g48641 not n18278 ; n18278_not
g48642 not n19178 ; n19178_not
g48643 not n11789 ; n11789_not
g48644 not n19574 ; n19574_not
g48645 not n11798 ; n11798_not
g48646 not n24767 ; n24767_not
g48647 not n24677 ; n24677_not
g48648 not n19952 ; n19952_not
g48649 not n15587 ; n15587_not
g48650 not n19169 ; n19169_not
g48651 not n15929 ; n15929_not
g48652 not n11969 ; n11969_not
g48653 not n22679 ; n22679_not
g48654 not n19727 ; n19727_not
g48655 not n25991 ; n25991_not
g48656 not n21986 ; n21986_not
g48657 not n22688 ; n22688_not
g48658 not n24668 ; n24668_not
g48659 not n20879 ; n20879_not
g48660 not n17666 ; n17666_not
g48661 not n14678 ; n14678_not
g48662 not n15569 ; n15569_not
g48663 not n16199 ; n16199_not
g48664 not n26189 ; n26189_not
g48665 not n19664 ; n19664_not
g48666 not n17909 ; n17909_not
g48667 not n11987 ; n11987_not
g48668 not n26198 ; n26198_not
g48669 not n25559 ; n25559_not
g48670 not n17675 ; n17675_not
g48671 not n19754 ; n19754_not
g48672 not n23939 ; n23939_not
g48673 not n19475 ; n19475_not
g48674 not n20969 ; n20969_not
g48675 not n18872 ; n18872_not
g48676 not n18890 ; n18890_not
g48677 not n14669 ; n14669_not
g48678 not n18629 ; n18629_not
g48679 not n18944 ; n18944_not
g48680 not n13967 ; n13967_not
g48681 not n16289 ; n16289_not
g48682 not n23876 ; n23876_not
g48683 not n20978 ; n20978_not
g48684 not n19763 ; n19763_not
g48685 not n18377 ; n18377_not
g48686 not n18638 ; n18638_not
g48687 not n18368 ; n18368_not
g48688 not n15983 ; n15983_not
g48689 not n24794 ; n24794_not
g48690 not n15866 ; n15866_not
g48691 not n22697 ; n22697_not
g48692 not n25586 ; n25586_not
g48693 not n17963 ; n17963_not
g48694 not n20897 ; n20897_not
g48695 not n13949 ; n13949_not
g48696 not n15578 ; n15578_not
g48697 not n19097 ; n19097_not
g48698 not n25577 ; n25577_not
g48699 not n17495 ; n17495_not
g48700 not n23498 ; n23498_not
g48701 not n15785 ; n15785_not
g48702 not n19088 ; n19088_not
g48703 not n17486 ; n17486_not
g48704 not n19079 ; n19079_not
g48705 not n13958 ; n13958_not
g48706 not n18980 ; n18980_not
g48707 not n21689 ; n21689_not
g48708 not n25568 ; n25568_not
g48709 not n19268 ; n19268_not
g48710 not n25694 ; n25694_not
g48711 not n19691 ; n19691_not
g48712 not n17972 ; n17972_not
g48713 not n23399 ; n23399_not
g48714 not n22598 ; n22598_not
g48715 not n15758 ; n15758_not
g48716 not n11879 ; n11879_not
g48717 not n11897 ; n11897_not
g48718 not n11888 ; n11888_not
g48719 not n25649 ; n25649_not
g48720 not n25685 ; n25685_not
g48721 not n20798 ; n20798_not
g48722 not n18566 ; n18566_not
g48723 not n23885 ; n23885_not
g48724 not n15668 ; n15668_not
g48725 not n17585 ; n17585_not
g48726 not n15749 ; n15749_not
g48727 not n13886 ; n13886_not
g48728 not n25829 ; n25829_not
g48729 not n25676 ; n25676_not
g48730 not n15776 ; n15776_not
g48731 not n15659 ; n15659_not
g48732 not n14768 ; n14768_not
g48733 not n25667 ; n25667_not
g48734 not n25793 ; n25793_not
g48735 not n25739 ; n25739_not
g48736 not n23777 ; n23777_not
g48737 not n18557 ; n18557_not
g48738 not n15695 ; n15695_not
g48739 not n24749 ; n24749_not
g48740 not n25748 ; n25748_not
g48741 not n19682 ; n19682_not
g48742 not n14786 ; n14786_not
g48743 not n23894 ; n23894_not
g48744 not n19385 ; n19385_not
g48745 not n19259 ; n19259_not
g48746 not n25757 ; n25757_not
g48747 not n15686 ; n15686_not
g48748 not n25766 ; n25766_not
g48749 not n17594 ; n17594_not
g48750 not n20789 ; n20789_not
g48751 not n24758 ; n24758_not
g48752 not n22499 ; n22499_not
g48753 not n23966 ; n23966_not
g48754 not n15677 ; n15677_not
g48755 not n25784 ; n25784_not
g48756 not n19934 ; n19934_not
g48757 not n15857 ; n15857_not
g48758 not n19196 ; n19196_not
g48759 not n17549 ; n17549_not
g48760 not n24695 ; n24695_not
g48761 not n19187 ; n19187_not
g48762 not n15875 ; n15875_not
g48763 not n25946 ; n25946_not
g48764 not n25937 ; n25937_not
g48765 not n18359 ; n18359_not
g48766 not n19718 ; n19718_not
g48767 not n24776 ; n24776_not
g48768 not n15884 ; n15884_not
g48769 not n25964 ; n25964_not
g48770 not n17657 ; n17657_not
g48771 not n25973 ; n25973_not
g48772 not n25982 ; n25982_not
g48773 not n15596 ; n15596_not
g48774 not n13877 ; n13877_not
g48775 not n25838 ; n25838_not
g48776 not n12788 ; n12788_not
g48777 not n25847 ; n25847_not
g48778 not n15794 ; n15794_not
g48779 not n18449 ; n18449_not
g48780 not n25856 ; n25856_not
g48781 not n18575 ; n18575_not
g48782 not n25865 ; n25865_not
g48783 not n17576 ; n17576_not
g48784 not n19277 ; n19277_not
g48785 not n17567 ; n17567_not
g48786 not n17981 ; n17981_not
g48787 not n25874 ; n25874_not
g48788 not n15839 ; n15839_not
g48789 not n25883 ; n25883_not
g48790 not n17558 ; n17558_not
g48791 not n19943 ; n19943_not
g48792 not n15848 ; n15848_not
g48793 not n25919 ; n25919_not
g48794 not n19844 ; n19844_not
g48795 not n16784 ; n16784_not
g48796 not n26855 ; n26855_not
g48797 not n23669 ; n23669_not
g48798 not n18665 ; n18665_not
g48799 not n13679 ; n13679_not
g48800 not n26828 ; n26828_not
g48801 not n16775 ; n16775_not
g48802 not n26837 ; n26837_not
g48803 not n16766 ; n16766_not
g48804 not n18467 ; n18467_not
g48805 not n17099 ; n17099_not
g48806 not n16757 ; n16757_not
g48807 not n18197 ; n18197_not
g48808 not n26945 ; n26945_not
g48809 not n23795 ; n23795_not
g48810 not n16829 ; n16829_not
g48811 not n26891 ; n26891_not
g48812 not n19853 ; n19853_not
g48813 not n18782 ; n18782_not
g48814 not n26927 ; n26927_not
g48815 not n26918 ; n26918_not
g48816 not n13589 ; n13589_not
g48817 not n23678 ; n23678_not
g48818 not n26909 ; n26909_not
g48819 not n18809 ; n18809_not
g48820 not n26882 ; n26882_not
g48821 not n26873 ; n26873_not
g48822 not n26729 ; n26729_not
g48823 not n26756 ; n26756_not
g48824 not n17198 ; n17198_not
g48825 not n16694 ; n16694_not
g48826 not n18179 ; n18179_not
g48827 not n26747 ; n26747_not
g48828 not n16685 ; n16685_not
g48829 not n18773 ; n18773_not
g48830 not n24479 ; n24479_not
g48831 not n26738 ; n26738_not
g48832 not n19826 ; n19826_not
g48833 not n13688 ; n13688_not
g48834 not n23975 ; n23975_not
g48835 not n16667 ; n16667_not
g48836 not n26819 ; n26819_not
g48837 not n18188 ; n18188_not
g48838 not n23984 ; n23984_not
g48839 not n16739 ; n16739_not
g48840 not n18827 ; n18827_not
g48841 not n18818 ; n18818_not
g48842 not n26792 ; n26792_not
g48843 not n26783 ; n26783_not
g48844 not n19835 ; n19835_not
g48845 not n17189 ; n17189_not
g48846 not n27197 ; n27197_not
g48847 not n13976 ; n13976_not
g48848 not n18395 ; n18395_not
g48849 not n16982 ; n16982_not
g48850 not n16919 ; n16919_not
g48851 not n24398 ; n24398_not
g48852 not n27188 ; n27188_not
g48853 not n18719 ; n18719_not
g48854 not n23993 ; n23993_not
g48855 not n27179 ; n27179_not
g48856 not n16856 ; n16856_not
g48857 not n18683 ; n18683_not
g48858 not n18728 ; n18728_not
g48859 not n27296 ; n27296_not
g48860 not n16964 ; n16964_not
g48861 not n18692 ; n18692_not
g48862 not n27287 ; n27287_not
g48863 not n18269 ; n18269_not
g48864 not n19871 ; n19871_not
g48865 not n27278 ; n27278_not
g48866 not n27269 ; n27269_not
g48867 not n16973 ; n16973_not
g48868 not n16946 ; n16946_not
g48869 not n16937 ; n16937_not
g48870 not n24389 ; n24389_not
g48871 not n14489 ; n14489_not
g48872 not n14498 ; n14498_not
g48873 not n18674 ; n18674_not
g48874 not n26990 ; n26990_not
g48875 not n26981 ; n26981_not
g48876 not n18791 ; n18791_not
g48877 not n16847 ; n16847_not
g48878 not n26972 ; n26972_not
g48879 not n16838 ; n16838_not
g48880 not n26963 ; n26963_not
g48881 not n13598 ; n13598_not
g48882 not n23687 ; n23687_not
g48883 not n26936 ; n26936_not
g48884 not n26954 ; n26954_not
g48885 not n16883 ; n16883_not
g48886 not n18737 ; n18737_not
g48887 not n27098 ; n27098_not
g48888 not n27089 ; n27089_not
g48889 not n16874 ; n16874_not
g48890 not n18746 ; n18746_not
g48891 not n19862 ; n19862_not
g48892 not n18755 ; n18755_not
g48893 not n23696 ; n23696_not
g48894 not n18764 ; n18764_not
g48895 not n16478 ; n16478_not
g48896 not n17387 ; n17387_not
g48897 not n18953 ; n18953_not
g48898 not n23957 ; n23957_not
g48899 not n19772 ; n19772_not
g48900 not n26396 ; n26396_not
g48901 not n17396 ; n17396_not
g48902 not n18962 ; n18962_not
g48903 not n26378 ; n26378_not
g48904 not n24569 ; n24569_not
g48905 not n21959 ; n21959_not
g48906 not n26369 ; n26369_not
g48907 not n10898 ; n10898_not
g48908 not n24578 ; n24578_not
g48909 not n18926 ; n18926_not
g48910 not n19790 ; n19790_not
g48911 not n26468 ; n26468_not
g48912 not n13994 ; n13994_not
g48913 not n26459 ; n26459_not
g48914 not n21896 ; n21896_not
g48915 not n21887 ; n21887_not
g48916 not n19781 ; n19781_not
g48917 not n18935 ; n18935_not
g48918 not n17369 ; n17369_not
g48919 not n16487 ; n16487_not
g48920 not n18098 ; n18098_not
g48921 not n17378 ; n17378_not
g48922 not n23948 ; n23948_not
g48923 not n17459 ; n17459_not
g48924 not n10988 ; n10988_not
g48925 not n18656 ; n18656_not
g48926 not n16379 ; n16379_not
g48927 not n10997 ; n10997_not
g48928 not n24596 ; n24596_not
g48929 not n20996 ; n20996_not
g48930 not n17468 ; n17468_not
g48931 not n21968 ; n21968_not
g48932 not n18647 ; n18647_not
g48933 not n20987 ; n20987_not
g48934 not n19970 ; n19970_not
g48935 not n18971 ; n18971_not
g48936 not n18089 ; n18089_not
g48937 not n21977 ; n21977_not
g48938 not n21788 ; n21788_not
g48939 not n13985 ; n13985_not
g48940 not n24587 ; n24587_not
g48941 not n10979 ; n10979_not
g48942 not n26297 ; n26297_not
g48943 not n16397 ; n16397_not
g48944 not n26288 ; n26288_not
g48945 not n17837 ; n17837_not
g48946 not n23759 ; n23759_not
g48947 not n26648 ; n26648_not
g48948 not n23849 ; n23849_not
g48949 not n18863 ; n18863_not
g48950 not n26639 ; n26639_not
g48951 not n19880 ; n19880_not
g48952 not n19817 ; n19817_not
g48953 not n16595 ; n16595_not
g48954 not n16586 ; n16586_not
g48955 not n18881 ; n18881_not
g48956 not n13499 ; n13499_not
g48957 not n26594 ; n26594_not
g48958 not n26576 ; n26576_not
g48959 not n18854 ; n18854_not
g48960 not n24488 ; n24488_not
g48961 not n21698 ; n21698_not
g48962 not n26693 ; n26693_not
g48963 not n16955 ; n16955_not
g48964 not n26684 ; n26684_not
g48965 not n16658 ; n16658_not
g48966 not n26675 ; n26675_not
g48967 not n14588 ; n14588_not
g48968 not n16649 ; n16649_not
g48969 not n26666 ; n26666_not
g48970 not n26657 ; n26657_not
g48971 not n16892 ; n16892_not
g48972 not n16568 ; n16568_not
g48973 not n23588 ; n23588_not
g48974 not n16559 ; n16559_not
g48975 not n18908 ; n18908_not
g48976 not n17297 ; n17297_not
g48977 not n20888 ; n20888_not
g48978 not n18917 ; n18917_not
g48979 not n18386 ; n18386_not
g48980 not n21869 ; n21869_not
g48981 not n26486 ; n26486_not
g48982 not n26477 ; n26477_not
g48983 not n21878 ; n21878_not
g48984 not n16496 ; n16496_not
g48985 not n23597 ; n23597_not
g48986 not n21779 ; n21779_not
g48987 not n16577 ; n16577_not
g48988 not n17279 ; n17279_not
g48989 not n13868 ; n13868_not
g48990 not n19808 ; n19808_not
g48991 not n26558 ; n26558_not
g48992 not n21797 ; n21797_not
g48993 not n13697 ; n13697_not
g48994 not n26549 ; n26549_not
g48995 not n19745 ; n19745_not
g48996 not n24947 ; n24947_not
g48997 not n14957 ; n14957_not
g48998 not n17882 ; n17882_not
g48999 not n19592 ; n19592_not
g49000 not n19565 ; n19565_not
g49001 not n24848 ; n24848_not
g49002 not n17918 ; n17918_not
g49003 not n17864 ; n17864_not
g49004 not n17738 ; n17738_not
g49005 not n14993 ; n14993_not
g49006 not n17783 ; n17783_not
g49007 not n19493 ; n19493_not
g49008 not n12779 ; n12779_not
g49009 not n13778 ; n13778_not
g49010 not n25199 ; n25199_not
g49011 not n25478 ; n25478_not
g49012 not n14876 ; n14876_not
g49013 not n12599 ; n12599_not
g49014 not n12959 ; n12959_not
g49015 not n24857 ; n24857_not
g49016 not n19457 ; n19457_not
g49017 not n24839 ; n24839_not
g49018 not n19358 ; n19358_not
g49019 not n15479 ; n15479_not
g49020 not n24992 ; n24992_not
g49021 not n19556 ; n19556_not
g49022 not n19925 ; n19925_not
g49023 not n14975 ; n14975_not
g49024 not n22949 ; n22949_not
g49025 not n22796 ; n22796_not
g49026 not n19439 ; n19439_not
g49027 not n19349 ; n19349_not
g49028 not n17747 ; n17747_not
g49029 not n18485 ; n18485_not
g49030 not n12869 ; n12869_not
g49031 not n19448 ; n19448_not
g49032 not n22886 ; n22886_not
g49033 not n14984 ; n14984_not
g49034 not n22958 ; n22958_not
g49035 not n12986 ; n12986_not
g49036 not n15497 ; n15497_not
g49037 not n24929 ; n24929_not
g49038 not n14399 ; n14399_not
g49039 not n12977 ; n12977_not
g49040 not n12968 ; n12968_not
g49041 not n19394 ; n19394_not
g49042 not n25298 ; n25298_not
g49043 not n17927 ; n17927_not
g49044 not n22994 ; n22994_not
g49045 not n14948 ; n14948_not
g49046 not n12797 ; n12797_not
g49047 not n22976 ; n22976_not
g49048 not n13769 ; n13769_not
g49049 not n18458 ; n18458_not
g49050 not n17756 ; n17756_not
g49051 not n22859 ; n22859_not
g49052 not n24884 ; n24884_not
g49053 not n19484 ; n19484_not
g49054 not n19583 ; n19583_not
g49055 not n13796 ; n13796_not
g49056 not n22868 ; n22868_not
g49057 not n17792 ; n17792_not
g49058 not n19619 ; n19619_not
g49059 not n17891 ; n17891_not
g49060 not n24938 ; n24938_not
g49061 not n14858 ; n14858_not
g49062 not n25469 ; n25469_not
g49063 not n17945 ; n17945_not
g49064 not n22877 ; n22877_not
g49065 not n25289 ; n25289_not
g49066 not n23858 ; n23858_not
g49067 not n19367 ; n19367_not
g49068 not n14966 ; n14966_not
g49069 not n14885 ; n14885_not
g49070 not n24956 ; n24956_not
g49071 not n24893 ; n24893_not
g49072 not n19466 ; n19466_not
g49073 not n19547 ; n19547_not
g49074 not n22778 ; n22778_not
g49075 not n19916 ; n19916_not
g49076 not n19673 ; n19673_not
g49077 not n11996 ; n11996_not
g49078 not n12689 ; n12689_not
g49079 not n23867 ; n23867_not
g49080 not n24983 ; n24983_not
g49081 not n12878 ; n12878_not
g49082 not n13859 ; n13859_not
g49083 not n12896 ; n12896_not
g49084 not n13787 ; n13787_not
g49085 not n22769 ; n22769_not
g49086 not n25388 ; n25388_not
g49087 not n18476 ; n18476_not
g49088 not n17774 ; n17774_not
g49089 not n14939 ; n14939_not
g49090 not n15389 ; n15389_not
g49091 not n17855 ; n17855_not
g49092 not n25397 ; n25397_not
g49093 not n22895 ; n22895_not
g49094 not n24974 ; n24974_not
g49095 not n19655 ; n19655_not
g49096 not n19529 ; n19529_not
g49097 not n25487 ; n25487_not
g49098 not n17828 ; n17828_not
g49099 not n15398 ; n15398_not
g49100 not n18494 ; n18494_not
g49101 not n15299 ; n15299_not
g49102 not n17936 ; n17936_not
g49103 not n24299 ; n24299_not
g49104 not n24875 ; n24875_not
g49105 not n22787 ; n22787_not
g49106 not n12698 ; n12698_not
g49107 not n25379 ; n25379_not
g49108 not n18539 ; n18539_not
g49109 not n19538 ; n19538_not
g49110 not n22967 ; n22967_not
g49111 not n17846 ; n17846_not
g49112 not n18296 ; n18296_not
g49113 not n19907 ; n19907_not
g49114 not n12887 ; n12887_not
g49115 not n17693 ; n17693_not
g49116 not n14894 ; n14894_not
g49117 not n17819 ; n17819_not
g49118 not n19637 ; n19637_not
g49119 not n14976 ; n14976_not
g49120 not n19089 ; n19089_not
g49121 not n26937 ; n26937_not
g49122 not n15768 ; n15768_not
g49123 not n13797 ; n13797_not
g49124 not n24687 ; n24687_not
g49125 not n14589 ; n14589_not
g49126 not n23985 ; n23985_not
g49127 not n15885 ; n15885_not
g49128 not n25983 ; n25983_not
g49129 not n25947 ; n25947_not
g49130 not n19476 ; n19476_not
g49131 not n18774 ; n18774_not
g49132 not n26199 ; n26199_not
g49133 not n19188 ; n19188_not
g49134 not n18792 ; n18792_not
g49135 not n15876 ; n15876_not
g49136 not n26766 ; n26766_not
g49137 not n19719 ; n19719_not
g49138 not n26946 ; n26946_not
g49139 not n22977 ; n22977_not
g49140 not n17388 ; n17388_not
g49141 not n19584 ; n19584_not
g49142 not n19854 ; n19854_not
g49143 not n25965 ; n25965_not
g49144 not n14679 ; n14679_not
g49145 not n17478 ; n17478_not
g49146 not n12888 ; n12888_not
g49147 not n17928 ; n17928_not
g49148 not n13959 ; n13959_not
g49149 not n19890 ; n19890_not
g49150 not n14688 ; n14688_not
g49151 not n25974 ; n25974_not
g49152 not n19467 ; n19467_not
g49153 not n23499 ; n23499_not
g49154 not n17487 ; n17487_not
g49155 not n19746 ; n19746_not
g49156 not n15966 ; n15966_not
g49157 not n15867 ; n15867_not
g49158 not n13779 ; n13779_not
g49159 not n16776 ; n16776_not
g49160 not n17676 ; n17676_not
g49161 not n18495 ; n18495_not
g49162 not n11799 ; n11799_not
g49163 not n14985 ; n14985_not
g49164 not n22869 ; n22869_not
g49165 not n26838 ; n26838_not
g49166 not n16767 ; n16767_not
g49167 not n15984 ; n15984_not
g49168 not n18585 ; n18585_not
g49169 not n19593 ; n19593_not
g49170 not n18198 ; n18198_not
g49171 not n19782 ; n19782_not
g49172 not n19179 ; n19179_not
g49173 not n22887 ; n22887_not
g49174 not n26865 ; n26865_not
g49175 not n16785 ; n16785_not
g49176 not n19728 ; n19728_not
g49177 not n15939 ; n15939_not
g49178 not n18387 ; n18387_not
g49179 not n24876 ; n24876_not
g49180 not n24669 ; n24669_not
g49181 not n19953 ; n19953_not
g49182 not n26856 ; n26856_not
g49183 not n17991 ; n17991_not
g49184 not n15948 ; n15948_not
g49185 not n18369 ; n18369_not
g49186 not n19449 ; n19449_not
g49187 not n26874 ; n26874_not
g49188 not n20799 ; n20799_not
g49189 not n19827 ; n19827_not
g49190 not n17919 ; n17919_not
g49191 not n18189 ; n18189_not
g49192 not n18468 ; n18468_not
g49193 not n18828 ; n18828_not
g49194 not n20898 ; n20898_not
g49195 not n19836 ; n19836_not
g49196 not n16578 ; n16578_not
g49197 not n19098 ; n19098_not
g49198 not n17496 ; n17496_not
g49199 not n19458 ; n19458_not
g49200 not n24948 ; n24948_not
g49201 not n26919 ; n26919_not
g49202 not n26784 ; n26784_not
g49203 not n26793 ; n26793_not
g49204 not n25992 ; n25992_not
g49205 not n26829 ; n26829_not
g49206 not n15993 ; n15993_not
g49207 not n12879 ; n12879_not
g49208 not n26892 ; n26892_not
g49209 not n25758 ; n25758_not
g49210 not n16758 ; n16758_not
g49211 not n18819 ; n18819_not
g49212 not n17775 ; n17775_not
g49213 not n17883 ; n17883_not
g49214 not n26739 ; n26739_not
g49215 not n24867 ; n24867_not
g49216 not n25875 ; n25875_not
g49217 not n14697 ; n14697_not
g49218 not n16749 ; n16749_not
g49219 not n15894 ; n15894_not
g49220 not n14994 ; n14994_not
g49221 not n18279 ; n18279_not
g49222 not n13788 ; n13788_not
g49223 not n26595 ; n26595_not
g49224 not n17856 ; n17856_not
g49225 not n18945 ; n18945_not
g49226 not n16479 ; n16479_not
g49227 not n23958 ; n23958_not
g49228 not n17379 ; n17379_not
g49229 not n23796 ; n23796_not
g49230 not n16488 ; n16488_not
g49231 not n26586 ; n26586_not
g49232 not n18936 ; n18936_not
g49233 not n18099 ; n18099_not
g49234 not n19980 ; n19980_not
g49235 not n21897 ; n21897_not
g49236 not n26577 ; n26577_not
g49237 not n14886 ; n14886_not
g49238 not n23598 ; n23598_not
g49239 not n16938 ; n16938_not
g49240 not n12969 ; n12969_not
g49241 not n17937 ; n17937_not
g49242 not n26379 ; n26379_not
g49243 not n23967 ; n23967_not
g49244 not n16596 ; n16596_not
g49245 not n19818 ; n19818_not
g49246 not n18486 ; n18486_not
g49247 not n19773 ; n19773_not
g49248 not n18666 ; n18666_not
g49249 not n19557 ; n19557_not
g49250 not n18963 ; n18963_not
g49251 not n17397 ; n17397_not
g49252 not n26397 ; n26397_not
g49253 not n13698 ; n13698_not
g49254 not n16587 ; n16587_not
g49255 not n14598 ; n14598_not
g49256 not n18873 ; n18873_not
g49257 not n18747 ; n18747_not
g49258 not n18918 ; n18918_not
g49259 not n19638 ; n19638_not
g49260 not n21789 ; n21789_not
g49261 not n26559 ; n26559_not
g49262 not n19548 ; n19548_not
g49263 not n19881 ; n19881_not
g49264 not n16983 ; n16983_not
g49265 not n18891 ; n18891_not
g49266 not n21798 ; n21798_not
g49267 not n17298 ; n17298_not
g49268 not n18909 ; n18909_not
g49269 not n19539 ; n19539_not
g49270 not n19917 ; n19917_not
g49271 not n23589 ; n23589_not
g49272 not n16569 ; n16569_not
g49273 not n17289 ; n17289_not
g49274 not n21888 ; n21888_not
g49275 not n14895 ; n14895_not
g49276 not n18576 ; n18576_not
g49277 not n17829 ; n17829_not
g49278 not n18927 ; n18927_not
g49279 not n19791 ; n19791_not
g49280 not n26469 ; n26469_not
g49281 not n18477 ; n18477_not
g49282 not n17847 ; n17847_not
g49283 not n21879 ; n21879_not
g49284 not n19809 ; n19809_not
g49285 not n22968 ; n22968_not
g49286 not n26568 ; n26568_not
g49287 not n19971 ; n19971_not
g49288 not n26487 ; n26487_not
g49289 not n26496 ; n26496_not
g49290 not n17748 ; n17748_not
g49291 not n12699 ; n12699_not
g49292 not n20889 ; n20889_not
g49293 not n24894 ; n24894_not
g49294 not n12789 ; n12789_not
g49295 not n21969 ; n21969_not
g49296 not n23976 ; n23976_not
g49297 not n18648 ; n18648_not
g49298 not n10989 ; n10989_not
g49299 not n23949 ; n23949_not
g49300 not n10998 ; n10998_not
g49301 not n19485 ; n19485_not
g49302 not n24597 ; n24597_not
g49303 not n24885 ; n24885_not
g49304 not n20988 ; n20988_not
g49305 not n18657 ; n18657_not
g49306 not n17199 ; n17199_not
g49307 not n16668 ; n16668_not
g49308 not n17874 ; n17874_not
g49309 not n17973 ; n17973_not
g49310 not n16389 ; n16389_not
g49311 not n26289 ; n26289_not
g49312 not n17793 ; n17793_not
g49313 not n19755 ; n19755_not
g49314 not n13689 ; n13689_not
g49315 not n26658 ; n26658_not
g49316 not n17469 ; n17469_not
g49317 not n26748 ; n26748_not
g49318 not n19575 ; n19575_not
g49319 not n16686 ; n16686_not
g49320 not n12798 ; n12798_not
g49321 not n13968 ; n13968_not
g49322 not n20979 ; n20979_not
g49323 not n26694 ; n26694_not
g49324 not n22995 ; n22995_not
g49325 not n25299 ; n25299_not
g49326 not n18639 ; n18639_not
g49327 not n19764 ; n19764_not
g49328 not n18837 ; n18837_not
g49329 not n21987 ; n21987_not
g49330 not n18981 ; n18981_not
g49331 not n26298 ; n26298_not
g49332 not n13986 ; n13986_not
g49333 not n12978 ; n12978_not
g49334 not n21978 ; n21978_not
g49335 not n24579 ; n24579_not
g49336 not n18972 ; n18972_not
g49337 not n26649 ; n26649_not
g49338 not n13977 ; n13977_not
g49339 not n14769 ; n14769_not
g49340 not n10899 ; n10899_not
g49341 not n14787 ; n14787_not
g49342 not n18864 ; n18864_not
g49343 not n16398 ; n16398_not
g49344 not n14877 ; n14877_not
g49345 not n24984 ; n24984_not
g49346 not n18855 ; n18855_not
g49347 not n24489 ; n24489_not
g49348 not n21699 ; n21699_not
g49349 not n24588 ; n24588_not
g49350 not n17784 ; n17784_not
g49351 not n26685 ; n26685_not
g49352 not n17865 ; n17865_not
g49353 not n19566 ; n19566_not
g49354 not n18990 ; n18990_not
g49355 not n26667 ; n26667_not
g49356 not n21996 ; n21996_not
g49357 not n19494 ; n19494_not
g49358 not n24498 ; n24498_not
g49359 not n18378 ; n18378_not
g49360 not n25749 ; n25749_not
g49361 not n16884 ; n16884_not
g49362 not n19683 ; n19683_not
g49363 not n19926 ; n19926_not
g49364 not n17586 ; n17586_not
g49365 not n19368 ; n19368_not
g49366 not n24957 ; n24957_not
g49367 not n25767 ; n25767_not
g49368 not n16875 ; n16875_not
g49369 not n25776 ; n25776_not
g49370 not n19863 ; n19863_not
g49371 not n25785 ; n25785_not
g49372 not n23697 ; n23697_not
g49373 not n24849 ; n24849_not
g49374 not n18549 ; n18549_not
g49375 not n16866 ; n16866_not
g49376 not n11898 ; n11898_not
g49377 not n17739 ; n17739_not
g49378 not n19359 ; n19359_not
g49379 not n16893 ; n16893_not
g49380 not n18729 ; n18729_not
g49381 not n25479 ; n25479_not
g49382 not n19674 ; n19674_not
g49383 not n15687 ; n15687_not
g49384 not n25398 ; n25398_not
g49385 not n13887 ; n13887_not
g49386 not n17595 ; n17595_not
g49387 not n17946 ; n17946_not
g49388 not n18738 ; n18738_not
g49389 not n15696 ; n15696_not
g49390 not n23859 ; n23859_not
g49391 not n25596 ; n25596_not
g49392 not n27099 ; n27099_not
g49393 not n18558 ; n18558_not
g49394 not n15777 ; n15777_not
g49395 not n25794 ; n25794_not
g49396 not n14967 ; n14967_not
g49397 not n19386 ; n19386_not
g49398 not n25839 ; n25839_not
g49399 not n15786 ; n15786_not
g49400 not n19656 ; n19656_not
g49401 not n24858 ; n24858_not
g49402 not n15795 ; n15795_not
g49403 not n18783 ; n18783_not
g49404 not n19395 ; n19395_not
g49405 not n25857 ; n25857_not
g49406 not n18675 ; n18675_not
g49407 not n16848 ; n16848_not
g49408 not n17577 ; n17577_not
g49409 not n11889 ; n11889_not
g49410 not n18756 ; n18756_not
g49411 not n13896 ; n13896_not
g49412 not n14778 ; n14778_not
g49413 not n17757 ; n17757_not
g49414 not n18567 ; n18567_not
g49415 not n17955 ; n17955_not
g49416 not n18297 ; n18297_not
g49417 not n16857 ; n16857_not
g49418 not n17568 ; n17568_not
g49419 not n19278 ; n19278_not
g49420 not n18765 ; n18765_not
g49421 not n22878 ; n22878_not
g49422 not n11979 ; n11979_not
g49423 not n27288 ; n27288_not
g49424 not n19872 ; n19872_not
g49425 not n19935 ; n19935_not
g49426 not n16956 ; n16956_not
g49427 not n13869 ; n13869_not
g49428 not n27279 ; n27279_not
g49429 not n14796 ; n14796_not
g49430 not n19296 ; n19296_not
g49431 not n16947 ; n16947_not
g49432 not n24786 ; n24786_not
g49433 not n22779 ; n22779_not
g49434 not n15588 ; n15588_not
g49435 not n24777 ; n24777_not
g49436 not n16974 ; n16974_not
g49437 not n19665 ; n19665_not
g49438 not n23877 ; n23877_not
g49439 not n24696 ; n24696_not
g49440 not n19629 ; n19629_not
g49441 not n18693 ; n18693_not
g49442 not n16965 ; n16965_not
g49443 not n25569 ; n25569_not
g49444 not n27297 ; n27297_not
g49445 not n15579 ; n15579_not
g49446 not n22698 ; n22698_not
g49447 not n11997 ; n11997_not
g49448 not n25587 ; n25587_not
g49449 not n24975 ; n24975_not
g49450 not n24795 ; n24795_not
g49451 not n24768 ; n24768_not
g49452 not n24399 ; n24399_not
g49453 not n14949 ; n14949_not
g49454 not n17964 ; n17964_not
g49455 not n15669 ; n15669_not
g49456 not n15498 ; n15498_not
g49457 not n22599 ; n22599_not
g49458 not n18684 ; n18684_not
g49459 not n23778 ; n23778_not
g49460 not n25686 ; n25686_not
g49461 not n25488 ; n25488_not
g49462 not n25695 ; n25695_not
g49463 not n23886 ; n23886_not
g49464 not n17892 ; n17892_not
g49465 not n15678 ; n15678_not
g49466 not n14958 ; n14958_not
g49467 not n19269 ; n19269_not
g49468 not n15597 ; n15597_not
g49469 not n22788 ; n22788_not
g49470 not n17658 ; n17658_not
g49471 not n13878 ; n13878_not
g49472 not n24993 ; n24993_not
g49473 not n23868 ; n23868_not
g49474 not n17649 ; n17649_not
g49475 not n22797 ; n22797_not
g49476 not n25497 ; n25497_not
g49477 not n25668 ; n25668_not
g49478 not n27189 ; n27189_not
g49479 not n15849 ; n15849_not
g49480 not n23688 ; n23688_not
g49481 not n19197 ; n19197_not
g49482 not n23679 ; n23679_not
g49483 not n26973 ; n26973_not
g49484 not n18288 ; n18288_not
g49485 not n17766 ; n17766_not
g49486 not n25884 ; n25884_not
g49487 not n16839 ; n16839_not
g49488 not n25938 ; n25938_not
g49489 not n22896 ; n22896_not
g49490 not n17982 ; n17982_not
g49491 not n17559 ; n17559_not
g49492 not n12897 ; n12897_not
g49493 not n26991 ; n26991_not
g49494 not n26982 ; n26982_not
g49495 not n19908 ; n19908_not
g49496 not n15858 ; n15858_not
g49497 not n19944 ; n19944_not
g49498 not n15399 ; n15399_not
g49499 not n14859 ; n14859_not
g49500 not n26955 ; n26955_not
g49501 not n23994 ; n23994_not
g49502 not n25866 ; n25866_not
g49503 not n17965 ; n17965_not
g49504 not n19819 ; n19819_not
g49505 not n25498 ; n25498_not
g49506 not n26965 ; n26965_not
g49507 not n14797 ; n14797_not
g49508 not n24967 ; n24967_not
g49509 not n17398 ; n17398_not
g49510 not n18955 ; n18955_not
g49511 not n24868 ; n24868_not
g49512 not n23968 ; n23968_not
g49513 not n14599 ; n14599_not
g49514 not n17767 ; n17767_not
g49515 not n22897 ; n22897_not
g49516 not n19459 ; n19459_not
g49517 not n19873 ; n19873_not
g49518 not n19279 ; n19279_not
g49519 not n19558 ; n19558_not
g49520 not n26398 ; n26398_not
g49521 not n24994 ; n24994_not
g49522 not n17857 ; n17857_not
g49523 not n19990 ; n19990_not
g49524 not n19882 ; n19882_not
g49525 not n16588 ; n16588_not
g49526 not n25993 ; n25993_not
g49527 not n12898 ; n12898_not
g49528 not n26389 ; n26389_not
g49529 not n22798 ; n22798_not
g49530 not n23779 ; n23779_not
g49531 not n18685 ; n18685_not
g49532 not n18577 ; n18577_not
g49533 not n17893 ; n17893_not
g49534 not n26857 ; n26857_not
g49535 not n25669 ; n25669_not
g49536 not n15679 ; n15679_not
g49537 not n13996 ; n13996_not
g49538 not n21997 ; n21997_not
g49539 not n19945 ; n19945_not
g49540 not n26668 ; n26668_not
g49541 not n17947 ; n17947_not
g49542 not n24679 ; n24679_not
g49543 not n18991 ; n18991_not
g49544 not n19936 ; n19936_not
g49545 not n16993 ; n16993_not
g49546 not n15868 ; n15868_not
g49547 not n26677 ; n26677_not
g49548 not n16939 ; n16939_not
g49549 not n26686 ; n26686_not
g49550 not n16894 ; n16894_not
g49551 not n14788 ; n14788_not
g49552 not n15967 ; n15967_not
g49553 not n17866 ; n17866_not
g49554 not n17776 ; n17776_not
g49555 not n24589 ; n24589_not
g49556 not n15688 ; n15688_not
g49557 not n16399 ; n16399_not
g49558 not n26299 ; n26299_not
g49559 not n16876 ; n16876_not
g49560 not n26875 ; n26875_not
g49561 not n19657 ; n19657_not
g49562 not n18487 ; n18487_not
g49563 not n15895 ; n15895_not
g49564 not n16795 ; n16795_not
g49565 not n17974 ; n17974_not
g49566 not n24499 ; n24499_not
g49567 not n18973 ; n18973_not
g49568 not n25489 ; n25489_not
g49569 not n25687 ; n25687_not
g49570 not n14896 ; n14896_not
g49571 not n21979 ; n21979_not
g49572 not n26893 ; n26893_not
g49573 not n13987 ; n13987_not
g49574 not n16984 ; n16984_not
g49575 not n19909 ; n19909_not
g49576 not n18676 ; n18676_not
g49577 not n26659 ; n26659_not
g49578 not n19675 ; n19675_not
g49579 not n18856 ; n18856_not
g49580 not n18982 ; n18982_not
g49581 not n19495 ; n19495_not
g49582 not n21988 ; n21988_not
g49583 not n19918 ; n19918_not
g49584 not n23887 ; n23887_not
g49585 not n14869 ; n14869_not
g49586 not n19846 ; n19846_not
g49587 not n18694 ; n18694_not
g49588 not n27289 ; n27289_not
g49589 not n19648 ; n19648_not
g49590 not n25588 ; n25588_not
g49591 not n11998 ; n11998_not
g49592 not n26497 ; n26497_not
g49593 not n19189 ; n19189_not
g49594 not n16498 ; n16498_not
g49595 not n19639 ; n19639_not
g49596 not n23959 ; n23959_not
g49597 not n26488 ; n26488_not
g49598 not n18793 ; n18793_not
g49599 not n12979 ; n12979_not
g49600 not n24976 ; n24976_not
g49601 not n26956 ; n26956_not
g49602 not n26938 ; n26938_not
g49603 not n13879 ; n13879_not
g49604 not n26479 ; n26479_not
g49605 not n25939 ; n25939_not
g49606 not n26569 ; n26569_not
g49607 not n25597 ; n25597_not
g49608 not n19783 ; n19783_not
g49609 not n17848 ; n17848_not
g49610 not n19792 ; n19792_not
g49611 not n25948 ; n25948_not
g49612 not a[10] ; a[10]_not
g49613 not n17677 ; n17677_not
g49614 not n17929 ; n17929_not
g49615 not n19756 ; n19756_not
g49616 not n23878 ; n23878_not
g49617 not n18892 ; n18892_not
g49618 not n17839 ; n17839_not
g49619 not n27298 ; n27298_not
g49620 not n17299 ; n17299_not
g49621 not n19666 ; n19666_not
g49622 not n25957 ; n25957_not
g49623 not n23995 ; n23995_not
g49624 not n26947 ; n26947_not
g49625 not n17956 ; n17956_not
g49626 not n15877 ; n15877_not
g49627 not n19855 ; n19855_not
g49628 not n17686 ; n17686_not
g49629 not n19549 ; n19549_not
g49630 not n22996 ; n22996_not
g49631 not n18748 ; n18748_not
g49632 not n22699 ; n22699_not
g49633 not n18919 ; n18919_not
g49634 not n26587 ; n26587_not
g49635 not n17659 ; n17659_not
g49636 not n15859 ; n15859_not
g49637 not n13789 ; n13789_not
g49638 not n23797 ; n23797_not
g49639 not n25984 ; n25984_not
g49640 not n16579 ; n16579_not
g49641 not n17695 ; n17695_not
g49642 not n18928 ; n18928_not
g49643 not n24778 ; n24778_not
g49644 not n24985 ; n24985_not
g49645 not n15886 ; n15886_not
g49646 not n14977 ; n14977_not
g49647 not n18946 ; n18946_not
g49648 not n15598 ; n15598_not
g49649 not n23599 ; n23599_not
g49650 not n27199 ; n27199_not
g49651 not n15589 ; n15589_not
g49652 not n17389 ; n17389_not
g49653 not n18874 ; n18874_not
g49654 not n25975 ; n25975_not
g49655 not n16957 ; n16957_not
g49656 not n25966 ; n25966_not
g49657 not n19297 ; n19297_not
g49658 not n21889 ; n21889_not
g49659 not n16966 ; n16966_not
g49660 not n12889 ; n12889_not
g49661 not n19954 ; n19954_not
g49662 not n16948 ; n16948_not
g49663 not n24796 ; n24796_not
g49664 not n24787 ; n24787_not
g49665 not n21898 ; n21898_not
g49666 not n26578 ; n26578_not
g49667 not n24949 ; n24949_not
g49668 not n24688 ; n24688_not
g49669 not n19981 ; n19981_not
g49670 not n18667 ; n18667_not
g49671 not n14887 ; n14887_not
g49672 not n23869 ; n23869_not
g49673 not n16489 ; n16489_not
g49674 not n18937 ; n18937_not
g49675 not n19288 ; n19288_not
g49676 not n24958 ; n24958_not
g49677 not n22978 ; n22978_not
g49678 not n18469 ; n18469_not
g49679 not n17758 ; n17758_not
g49680 not n15949 ; n15949_not
g49681 not n26767 ; n26767_not
g49682 not n18757 ; n18757_not
g49683 not n18298 ; n18298_not
g49684 not n14689 ; n14689_not
g49685 not n19468 ; n19468_not
g49686 not n25876 ; n25876_not
g49687 not n16858 ; n16858_not
g49688 not n15958 ; n15958_not
g49689 not n17488 ; n17488_not
g49690 not n26776 ; n26776_not
g49691 not n17938 ; n17938_not
g49692 not n19729 ; n19729_not
g49693 not n22888 ; n22888_not
g49694 not n26785 ; n26785_not
g49695 not n15778 ; n15778_not
g49696 not n15769 ; n15769_not
g49697 not n22969 ; n22969_not
g49698 not n19747 ; n19747_not
g49699 not n19378 ; n19378_not
g49700 not n25777 ; n25777_not
g49701 not n19864 ; n19864_not
g49702 not n24877 ; n24877_not
g49703 not n17884 ; n17884_not
g49704 not n18496 ; n18496_not
g49705 not n22987 ; n22987_not
g49706 not n14878 ; n14878_not
g49707 not n16687 ; n16687_not
g49708 not n19828 ; n19828_not
g49709 not n17983 ; n17983_not
g49710 not n24886 ; n24886_not
g49711 not n16867 ; n16867_not
g49712 not n26749 ; n26749_not
g49713 not n19576 ; n19576_not
g49714 not n18388 ; n18388_not
g49715 not n25795 ; n25795_not
g49716 not n14779 ; n14779_not
g49717 not n23986 ; n23986_not
g49718 not n16768 ; n16768_not
g49719 not n17479 ; n17479_not
g49720 not n13897 ; n13897_not
g49721 not n19567 ; n19567_not
g49722 not n25849 ; n25849_not
g49723 not n18775 ; n18775_not
g49724 not n16759 ; n16759_not
g49725 not n15976 ; n15976_not
g49726 not n18784 ; n18784_not
g49727 not n17578 ; n17578_not
g49728 not n15796 ; n15796_not
g49729 not n18595 ; n18595_not
g49730 not n15994 ; n15994_not
g49731 not n16849 ; n16849_not
g49732 not n13798 ; n13798_not
g49733 not n25858 ; n25858_not
g49734 not n19396 ; n19396_not
g49735 not n18586 ; n18586_not
g49736 not n15985 ; n15985_not
g49737 not n19594 ; n19594_not
g49738 not n19099 ; n19099_not
g49739 not n26992 ; n26992_not
g49740 not n19738 ; n19738_not
g49741 not n26794 ; n26794_not
g49742 not n26848 ; n26848_not
g49743 not n17497 ; n17497_not
g49744 not n26758 ; n26758_not
g49745 not n17569 ; n17569_not
g49746 not n16777 ; n16777_not
g49747 not n19963 ; n19963_not
g49748 not n17785 ; n17785_not
g49749 not n19891 ; n19891_not
g49750 not n18829 ; n18829_not
g49751 not n14995 ; n14995_not
g49752 not n19927 ; n19927_not
g49753 not n14968 ; n14968_not
g49754 not n19837 ; n19837_not
g49755 not n14698 ; n14698_not
g49756 not n15787 ; n15787_not
g49757 not n24859 ; n24859_not
g49758 not n19387 ; n19387_not
g49759 not n18838 ; n18838_not
g49760 not n17749 ; n17749_not
g49761 not n16678 ; n16678_not
g49762 not n16885 ; n16885_not
g49763 not n25894 ; n25894_not
g49764 not n26866 ; n26866_not
g49765 not n26974 ; n26974_not
g49766 not n18649 ; n18649_not
g49767 not n18379 ; n18379_not
g49768 not n24895 ; n24895_not
g49769 not n20989 ; n20989_not
g49770 not n19765 ; n19765_not
g49771 not n14959 ; n14959_not
g49772 not n17587 ; n17587_not
g49773 not n18289 ; n18289_not
g49774 not n19684 ; n19684_not
g49775 not n25885 ; n25885_not
g49776 not n13888 ; n13888_not
g49777 not n17794 ; n17794_not
g49778 not n17596 ; n17596_not
g49779 not n12988 ; n12988_not
g49780 not n17992 ; n17992_not
g49781 not n18739 ; n18739_not
g49782 not n13978 ; n13978_not
g49783 not n15697 ; n15697_not
g49784 not n16669 ; n16669_not
g49785 not n18847 ; n18847_not
g49786 not n17875 ; n17875_not
g49787 not n18658 ; n18658_not
g49788 not n12997 ; n12997_not
g49789 not n19486 ; n19486_not
g49790 not n24598 ; n24598_not
g49791 not n10999 ; n10999_not
g49792 not n26695 ; n26695_not
g49793 not n19369 ; n19369_not
g49794 not n25768 ; n25768_not
g49795 not n25759 ; n25759_not
g49796 not n23698 ; n23698_not
g49797 not n14978 ; n14978_not
g49798 not n26939 ; n26939_not
g49799 not n26678 ; n26678_not
g49800 not n26867 ; n26867_not
g49801 not n16994 ; n16994_not
g49802 not n26885 ; n26885_not
g49803 not n18848 ; n18848_not
g49804 not n19388 ; n19388_not
g49805 not n19865 ; n19865_not
g49806 not n19838 ; n19838_not
g49807 not n17894 ; n17894_not
g49808 not n26669 ; n26669_not
g49809 not n24878 ; n24878_not
g49810 not n14969 ; n14969_not
g49811 not n17876 ; n17876_not
g49812 not n16688 ; n16688_not
g49813 not n23798 ; n23798_not
g49814 not n16886 ; n16886_not
g49815 not n17489 ; n17489_not
g49816 not n18389 ; n18389_not
g49817 not n23699 ; n23699_not
g49818 not n19856 ; n19856_not
g49819 not n26858 ; n26858_not
g49820 not n24995 ; n24995_not
g49821 not n18398 ; n18398_not
g49822 not n26696 ; n26696_not
g49823 not n18668 ; n18668_not
g49824 not n19595 ; n19595_not
g49825 not n26993 ; n26993_not
g49826 not a[11] ; a[11]_not
g49827 not n17867 ; n17867_not
g49828 not n16895 ; n16895_not
g49829 not n16859 ; n16859_not
g49830 not b[10] ; b[10]_not
g49831 not n18893 ; n18893_not
g49832 not n17759 ; n17759_not
g49833 not n18785 ; n18785_not
g49834 not n27299 ; n27299_not
g49835 not n16589 ; n16589_not
g49836 not n16787 ; n16787_not
g49837 not n12899 ; n12899_not
g49838 not n24968 ; n24968_not
g49839 not n19892 ; n19892_not
g49840 not n19829 ; n19829_not
g49841 not n26876 ; n26876_not
g49842 not n17885 ; n17885_not
g49843 not n19847 ; n19847_not
g49844 not n23996 ; n23996_not
g49845 not n19559 ; n19559_not
g49846 not n18884 ; n18884_not
g49847 not a[20] ; a[20]_not
g49848 not n26588 ; n26588_not
g49849 not n16769 ; n16769_not
g49850 not n18299 ; n18299_not
g49851 not n18758 ; n18758_not
g49852 not n18686 ; n18686_not
g49853 not n26966 ; n26966_not
g49854 not n26984 ; n26984_not
g49855 not n16796 ; n16796_not
g49856 not n19577 ; n19577_not
g49857 not n16778 ; n16778_not
g49858 not n18677 ; n18677_not
g49859 not n16697 ; n16697_not
g49860 not n26777 ; n26777_not
g49861 not n18794 ; n18794_not
g49862 not n26759 ; n26759_not
g49863 not n14879 ; n14879_not
g49864 not n19982 ; n19982_not
g49865 not n16679 ; n16679_not
g49866 not n26894 ; n26894_not
g49867 not n18776 ; n18776_not
g49868 not n18857 ; n18857_not
g49869 not n26768 ; n26768_not
g49870 not n19883 ; n19883_not
g49871 not n26849 ; n26849_not
g49872 not n16958 ; n16958_not
g49873 not n16985 ; n16985_not
g49874 not n16868 ; n16868_not
g49875 not n26957 ; n26957_not
g49876 not n26795 ; n26795_not
g49877 not n23987 ; n23987_not
g49878 not n17858 ; n17858_not
g49879 not n18839 ; n18839_not
g49880 not n19874 ; n19874_not
g49881 not n23969 ; n23969_not
g49882 not n14897 ; n14897_not
g49883 not n18749 ; n18749_not
g49884 not n18875 ; n18875_not
g49885 not n16949 ; n16949_not
g49886 not n16967 ; n16967_not
g49887 not n26786 ; n26786_not
g49888 not n19991 ; n19991_not
g49889 not n14996 ; n14996_not
g49890 not n24977 ; n24977_not
g49891 not n26975 ; n26975_not
g49892 not n25985 ; n25985_not
g49893 not n21989 ; n21989_not
g49894 not n15959 ; n15959_not
g49895 not n19955 ; n19955_not
g49896 not n15968 ; n15968_not
g49897 not n15977 ; n15977_not
g49898 not n17948 ; n17948_not
g49899 not n19739 ; n19739_not
g49900 not n15986 ; n15986_not
g49901 not n13799 ; n13799_not
g49902 not n15995 ; n15995_not
g49903 not n18596 ; n18596_not
g49904 not n18587 ; n18587_not
g49905 not n25949 ; n25949_not
g49906 not n25958 ; n25958_not
g49907 not n15878 ; n15878_not
g49908 not n24689 ; n24689_not
g49909 not n25967 ; n25967_not
g49910 not n25976 ; n25976_not
g49911 not n24869 ; n24869_not
g49912 not n25994 ; n25994_not
g49913 not n15887 ; n15887_not
g49914 not n17939 ; n17939_not
g49915 not n19919 ; n19919_not
g49916 not n17777 ; n17777_not
g49917 not n17993 ; n17993_not
g49918 not n19766 ; n19766_not
g49919 not n20999 ; n20999_not
g49920 not n12989 ; n12989_not
g49921 not n22997 ; n22997_not
g49922 not n19487 ; n19487_not
g49923 not n24896 ; n24896_not
g49924 not n13979 ; n13979_not
g49925 not n18659 ; n18659_not
g49926 not n17795 ; n17795_not
g49927 not n18992 ; n18992_not
g49928 not n21998 ; n21998_not
g49929 not n17786 ; n17786_not
g49930 not n14699 ; n14699_not
g49931 not n17498 ; n17498_not
g49932 not n19964 ; n19964_not
g49933 not n19748 ; n19748_not
g49934 not n19469 ; n19469_not
g49935 not n24887 ; n24887_not
g49936 not n19478 ; n19478_not
g49937 not n22988 ; n22988_not
g49938 not n24779 ; n24779_not
g49939 not n15599 ; n15599_not
g49940 not n17966 ; n17966_not
g49941 not n22799 ; n22799_not
g49942 not n25499 ; n25499_not
g49943 not n25679 ; n25679_not
g49944 not n12998 ; n12998_not
g49945 not n25688 ; n25688_not
g49946 not n23888 ; n23888_not
g49947 not n19676 ; n19676_not
g49948 not n15689 ; n15689_not
g49949 not n19928 ; n19928_not
g49950 not n15698 ; n15698_not
g49951 not n17588 ; n17588_not
g49952 not n19298 ; n19298_not
g49953 not n23789 ; n23789_not
g49954 not n17678 ; n17678_not
g49955 not n23879 ; n23879_not
g49956 not n18983 ; n18983_not
g49957 not n19667 ; n19667_not
g49958 not n19658 ; n19658_not
g49959 not n17669 ; n17669_not
g49960 not n17687 ; n17687_not
g49961 not n25589 ; n25589_not
g49962 not n11999 ; n11999_not
g49963 not n25598 ; n25598_not
g49964 not n24788 ; n24788_not
g49965 not n19289 ; n19289_not
g49966 not n17696 ; n17696_not
g49967 not n25859 ; n25859_not
g49968 not n17975 ; n17975_not
g49969 not n19397 ; n19397_not
g49970 not n25877 ; n25877_not
g49971 not n22889 ; n22889_not
g49972 not n25886 ; n25886_not
g49973 not n17984 ; n17984_not
g49974 not n25895 ; n25895_not
g49975 not n22898 ; n22898_not
g49976 not n24698 ; n24698_not
g49977 not n18578 ; n18578_not
g49978 not n17768 ; n17768_not
g49979 not n19649 ; n19649_not
g49980 not n15869 ; n15869_not
g49981 not n13889 ; n13889_not
g49982 not n23897 ; n23897_not
g49983 not n19685 ; n19685_not
g49984 not n25778 ; n25778_not
g49985 not n19379 ; n19379_not
g49986 not n19694 ; n19694_not
g49987 not n25796 ; n25796_not
g49988 not n13898 ; n13898_not
g49989 not n15779 ; n15779_not
g49990 not n17579 ; n17579_not
g49991 not n15788 ; n15788_not
g49992 not n25769 ; n25769_not
g49993 not n15797 ; n15797_not
g49994 not n26498 ; n26498_not
g49995 not n26489 ; n26489_not
g49996 not n18947 ; n18947_not
g49997 not n16499 ; n16499_not
g49998 not n19757 ; n19757_not
g49999 not n19784 ; n19784_not
g50000 not n19973 ; n19973_not
g50001 not n18938 ; n18938_not
g50002 not n14888 ; n14888_not
g50003 not n18956 ; n18956_not
g50004 not n19775 ; n19775_not
g50005 not n21899 ; n21899_not
g50006 not n18974 ; n18974_not
g50007 not n19793 ; n19793_not
g50008 not n22979 ; n22979_not
g50009 not n24797 ; n24797_not
g50010 not n13997 ; n13997_not
g50011 not n18488 ; n18488_not
g50012 not n13988 ; n13988_not
g50013 not n18929 ; n18929_not
g50014 not n17399 ; n17399_not
g50015 not n19884 ; n19884_not
g50016 not n19686 ; n19686_not
g50017 not n18885 ; n18885_not
g50018 not n18588 ; n18588_not
g50019 not n12999 ; n12999_not
g50020 not a[30] ; a[30]_not
g50021 not n17796 ; n17796_not
g50022 not n17499 ; n17499_not
g50023 not n15996 ; n15996_not
g50024 not n18966 ; n18966_not
g50025 not n24879 ; n24879_not
g50026 not n26976 ; n26976_not
g50027 not n13989 ; n13989_not
g50028 not a[21] ; a[21]_not
g50029 not n18759 ; n18759_not
g50030 not n25788 ; n25788_not
g50031 not n17589 ; n17589_not
g50032 not n14988 ; n14988_not
g50033 not n18948 ; n18948_not
g50034 not b[20] ; b[20]_not
g50035 not n26787 ; n26787_not
g50036 not n13998 ; n13998_not
g50037 not n16599 ; n16599_not
g50038 not n25896 ; n25896_not
g50039 not n25779 ; n25779_not
g50040 not n18399 ; n18399_not
g50041 not n18867 ; n18867_not
g50042 not n19857 ; n19857_not
g50043 not n19992 ; n19992_not
g50044 not n19893 ; n19893_not
g50045 not n17985 ; n17985_not
g50046 not n26967 ; n26967_not
g50047 not n17787 ; n17787_not
g50048 not n17859 ; n17859_not
g50049 not n19839 ; n19839_not
g50050 not n16977 ; n16977_not
g50051 not n17679 ; n17679_not
g50052 not n26589 ; n26589_not
g50053 not n26598 ; n26598_not
g50054 not n18597 ; n18597_not
g50055 not n24996 ; n24996_not
g50056 not n19794 ; n19794_not
g50057 not n18579 ; n18579_not
g50058 not n26796 ; n26796_not
g50059 not n24699 ; n24699_not
g50060 not n23889 ; n23889_not
g50061 not n19875 ; n19875_not
g50062 not n25599 ; n25599_not
g50063 not n26886 ; n26886_not
g50064 not n19938 ; n19938_not
g50065 not n18795 ; n18795_not
g50066 not n15879 ; n15879_not
g50067 not n25986 ; n25986_not
g50068 not n25878 ; n25878_not
g50069 not n16995 ; n16995_not
g50070 not n26895 ; n26895_not
g50071 not n15699 ; n15699_not
g50072 not n16896 ; n16896_not
g50073 not n16797 ; n16797_not
g50074 not n26859 ; n26859_not
g50075 not n25995 ; n25995_not
g50076 not n23988 ; n23988_not
g50077 not n16887 ; n16887_not
g50078 not n17598 ; n17598_not
g50079 not n16788 ; n16788_not
g50080 not n19929 ; n19929_not
g50081 not n26499 ; n26499_not
g50082 not n15888 ; n15888_not
g50083 not n15978 ; n15978_not
g50084 not n17769 ; n17769_not
g50085 not n15969 ; n15969_not
g50086 not n17967 ; n17967_not
g50087 not n16878 ; n16878_not
g50088 not n25689 ; n25689_not
g50089 not n19956 ; n19956_not
g50090 not n19596 ; n19596_not
g50091 not n16779 ; n16779_not
g50092 not n19983 ; n19983_not
g50093 not n25959 ; n25959_not
g50094 not n23799 ; n23799_not
g50095 not n25698 ; n25698_not
g50096 not n14979 ; n14979_not
g50097 not n17778 ; n17778_not
g50098 not n18876 ; n18876_not
g50099 not n25968 ; n25968_not
g50100 not n26868 ; n26868_not
g50101 not n19776 ; n19776_not
g50102 not n19848 ; n19848_not
g50103 not n25977 ; n25977_not
g50104 not n26877 ; n26877_not
g50105 not n19299 ; n19299_not
g50106 not n18975 ; n18975_not
g50107 not n18894 ; n18894_not
g50108 not n22998 ; n22998_not
g50109 not n18489 ; n18489_not
g50110 not n19767 ; n19767_not
g50111 not n17895 ; n17895_not
g50112 not n26679 ; n26679_not
g50113 not n19659 ; n19659_not
g50114 not n24978 ; n24978_not
g50115 not n17688 ; n17688_not
g50116 not n17958 ; n17958_not
g50117 not n19866 ; n19866_not
g50118 not n23979 ; n23979_not
g50119 not n25797 ; n25797_not
g50120 not n26994 ; n26994_not
g50121 not n17877 ; n17877_not
g50122 not n19758 ; n19758_not
g50123 not n22989 ; n22989_not
g50124 not n23898 ; n23898_not
g50125 not n16869 ; n16869_not
g50126 not n18669 ; n18669_not
g50127 not n19695 ; n19695_not
g50128 not n24798 ; n24798_not
g50129 not n18777 ; n18777_not
g50130 not n19488 ; n19488_not
g50131 not n26697 ; n26697_not
g50132 not n14799 ; n14799_not
g50133 not n19569 ; n19569_not
g50134 not n24969 ; n24969_not
g50135 not n18678 ; n18678_not
g50136 not n19389 ; n19389_not
g50137 not n19974 ; n19974_not
g50138 not n19497 ; n19497_not
g50139 not n24897 ; n24897_not
g50140 not n18849 ; n18849_not
g50141 not n16986 ; n16986_not
g50142 not a[12] ; a[12]_not
g50143 not n15798 ; n15798_not
g50144 not n16698 ; n16698_not
g50145 not n18939 ; n18939_not
g50146 not n21999 ; n21999_not
g50147 not n13899 ; n13899_not
g50148 not n19398 ; n19398_not
g50149 not n19578 ; n19578_not
g50150 not n17697 ; n17697_not
g50151 not n18858 ; n18858_not
g50152 not n19965 ; n19965_not
g50153 not n19668 ; n19668_not
g50154 not n26985 ; n26985_not
g50155 not n26769 ; n26769_not
g50156 not n18984 ; n18984_not
g50157 not n26778 ; n26778_not
g50158 not n18768 ; n18768_not
g50159 not n19587 ; n19587_not
g50160 not n24987 ; n24987_not
g50161 not n24789 ; n24789_not
g50162 not n16968 ; n16968_not
g50163 not n19785 ; n19785_not
g50164 not n14898 ; n14898_not
g50165 not b[11] ; b[11]_not
g50166 not n16689 ; n16689_not
g50167 not n18687 ; n18687_not
g50168 not n17976 ; n17976_not
g50169 not n24888 ; n24888_not
g50170 not n17868 ; n17868_not
g50171 not n17949 ; n17949_not
g50172 not n19479 ; n19479_not
g50173 not n25869 ; n25869_not
g50174 not n19786 ; n19786_not
g50175 not n18769 ; n18769_not
g50176 not n19597 ; n19597_not
g50177 not n18796 ; n18796_not
g50178 not n23989 ; n23989_not
g50179 not a[40] ; a[40]_not
g50180 not n18499 ; n18499_not
g50181 not n17977 ; n17977_not
g50182 not n25996 ; n25996_not
g50183 not n16987 ; n16987_not
g50184 not n26959 ; n26959_not
g50185 not n19696 ; n19696_not
g50186 not n18679 ; n18679_not
g50187 not n25987 ; n25987_not
g50188 not n26599 ; n26599_not
g50189 not n18886 ; n18886_not
g50190 not n16996 ; n16996_not
g50191 not n19687 ; n19687_not
g50192 not n17887 ; n17887_not
g50193 not n19867 ; n19867_not
g50194 not n19957 ; n19957_not
g50195 not n19948 ; n19948_not
g50196 not n26968 ; n26968_not
g50197 not n25897 ; n25897_not
g50198 not n26986 ; n26986_not
g50199 not n25879 ; n25879_not
g50200 not n19399 ; n19399_not
g50201 not n25789 ; n25789_not
g50202 not n26977 ; n26977_not
g50203 not n23899 ; n23899_not
g50204 not n25978 ; n25978_not
g50205 not n18778 ; n18778_not
g50206 not n25969 ; n25969_not
g50207 not n26878 ; n26878_not
g50208 not n17986 ; n17986_not
g50209 not n18877 ; n18877_not
g50210 not n18949 ; n18949_not
g50211 not n19795 ; n19795_not
g50212 not n17959 ; n17959_not
g50213 not n16879 ; n16879_not
g50214 not n15799 ; n15799_not
g50215 not n19858 ; n19858_not
g50216 not n26995 ; n26995_not
g50217 not n18688 ; n18688_not
g50218 not n19489 ; n19489_not
g50219 not n19993 ; n19993_not
g50220 not n16969 ; n16969_not
g50221 not n16699 ; n16699_not
g50222 not n19669 ; n19669_not
g50223 not n19579 ; n19579_not
g50224 not n19966 ; n19966_not
g50225 not n18859 ; n18859_not
g50226 not n24988 ; n24988_not
g50227 not n26779 ; n26779_not
g50228 not n19588 ; n19588_not
g50229 not b[21] ; b[21]_not
g50230 not n14998 ; n14998_not
g50231 not a[22] ; a[22]_not
g50232 not n19768 ; n19768_not
g50233 not n26797 ; n26797_not
g50234 not n17797 ; n17797_not
g50235 not n16978 ; n16978_not
g50236 not n18868 ; n18868_not
g50237 not n18589 ; n18589_not
g50238 not n18598 ; n18598_not
g50239 not n19876 ; n19876_not
g50240 not n18985 ; n18985_not
g50241 not n18976 ; n18976_not
g50242 not b[12] ; b[12]_not
g50243 not n19885 ; n19885_not
g50244 not n19498 ; n19498_not
g50245 not n18895 ; n18895_not
g50246 not a[13] ; a[13]_not
g50247 not n14899 ; n14899_not
g50248 not n26689 ; n26689_not
g50249 not n26698 ; n26698_not
g50250 not n24898 ; n24898_not
g50251 not n17869 ; n17869_not
g50252 not n24799 ; n24799_not
g50253 not n13999 ; n13999_not
g50254 not n18697 ; n18697_not
g50255 not n24979 ; n24979_not
g50256 not n17689 ; n17689_not
g50257 not n17878 ; n17878_not
g50258 not n19777 ; n19777_not
g50259 not n19759 ; n19759_not
g50260 not b[30] ; b[30]_not
g50261 not n17599 ; n17599_not
g50262 not n19984 ; n19984_not
g50263 not a[31] ; a[31]_not
g50264 not n17779 ; n17779_not
g50265 not n18958 ; n18958_not
g50266 not n25699 ; n25699_not
g50267 not n26869 ; n26869_not
g50268 not n15898 ; n15898_not
g50269 not n26896 ; n26896_not
g50270 not n25888 ; n25888_not
g50271 not n26887 ; n26887_not
g50272 not n19975 ; n19975_not
g50273 not n16789 ; n16789_not
g50274 not n24997 ; n24997_not
g50275 not n15997 ; n15997_not
g50276 not n16798 ; n16798_not
g50277 not n15889 ; n15889_not
g50278 not n18967 ; n18967_not
g50279 not n15988 ; n15988_not
g50280 not n17896 ; n17896_not
g50281 not n15979 ; n15979_not
g50282 not n14989 ; n14989_not
g50283 not b[31] ; b[31]_not
g50284 not b[40] ; b[40]_not
g50285 not a[23] ; a[23]_not
g50286 not n18986 ; n18986_not
g50287 not n19697 ; n19697_not
g50288 not a[32] ; a[32]_not
g50289 not n16889 ; n16889_not
g50290 not b[13] ; b[13]_not
g50291 not n19679 ; n19679_not
g50292 not n18896 ; n18896_not
g50293 not a[41] ; a[41]_not
g50294 not a[14] ; a[14]_not
g50295 not n24998 ; n24998_not
g50296 not n16979 ; n16979_not
g50297 not n17888 ; n17888_not
g50298 not b[22] ; b[22]_not
g50299 not a[50] ; a[50]_not
g50300 not n19886 ; n19886_not
g50301 not n19688 ; n19688_not
g50302 not n18698 ; n18698_not
g50303 not n17969 ; n17969_not
g50304 not n16988 ; n16988_not
g50305 not n19868 ; n19868_not
g50306 not n16997 ; n16997_not
g50307 not n17897 ; n17897_not
g50308 not n18689 ; n18689_not
g50309 not n19796 ; n19796_not
g50310 not n24989 ; n24989_not
g50311 not n18968 ; n18968_not
g50312 not n15989 ; n15989_not
g50313 not n18869 ; n18869_not
g50314 not n19985 ; n19985_not
g50315 not n19598 ; n19598_not
g50316 not n25979 ; n25979_not
g50317 not n17996 ; n17996_not
g50318 not n25997 ; n25997_not
g50319 not n26888 ; n26888_not
g50320 not n17987 ; n17987_not
g50321 not n15899 ; n15899_not
g50322 not n16799 ; n16799_not
g50323 not n18797 ; n18797_not
g50324 not n19778 ; n19778_not
g50325 not n25988 ; n25988_not
g50326 not n19949 ; n19949_not
g50327 not n23999 ; n23999_not
g50328 not n25898 ; n25898_not
g50329 not n25889 ; n25889_not
g50330 not n18995 ; n18995_not
g50331 not n19499 ; n19499_not
g50332 not n19769 ; n19769_not
g50333 not n18959 ; n18959_not
g50334 not n19877 ; n19877_not
g50335 not n19967 ; n19967_not
g50336 not n17879 ; n17879_not
g50337 not n19994 ; n19994_not
g50338 not n19589 ; n19589_not
g50339 not n14999 ; n14999_not
g50340 not n26798 ; n26798_not
g50341 not n19958 ; n19958_not
g50342 not n17798 ; n17798_not
g50343 not n15998 ; n15998_not
g50344 not n18599 ; n18599_not
g50345 not n18887 ; n18887_not
g50346 not n19895 ; n19895_not
g50347 not n18779 ; n18779_not
g50348 not n19859 ; n19859_not
g50349 not n18788 ; n18788_not
g50350 not n26996 ; n26996_not
g50351 not n26978 ; n26978_not
g50352 not b[23] ; b[23]_not
g50353 not a[51] ; a[51]_not
g50354 not a[60] ; a[60]_not
g50355 not n19896 ; n19896_not
g50356 not n18897 ; n18897_not
g50357 not b[50] ; b[50]_not
g50358 not a[24] ; a[24]_not
g50359 not n25998 ; n25998_not
g50360 not n26997 ; n26997_not
g50361 not a[15] ; a[15]_not
g50362 not n18969 ; n18969_not
g50363 not n18699 ; n18699_not
g50364 not n18798 ; n18798_not
g50365 not n19968 ; n19968_not
g50366 not n24999 ; n24999_not
g50367 not n25989 ; n25989_not
g50368 not b[41] ; b[41]_not
g50369 not a[42] ; a[42]_not
g50370 not n26898 ; n26898_not
g50371 not n17997 ; n17997_not
g50372 not n26799 ; n26799_not
g50373 not n19986 ; n19986_not
g50374 not n16989 ; n16989_not
g50375 not n17988 ; n17988_not
g50376 not n19689 ; n19689_not
g50377 not b[32] ; b[32]_not
g50378 not a[33] ; a[33]_not
g50379 not n26889 ; n26889_not
g50380 not n18789 ; n18789_not
g50381 not n19959 ; n19959_not
g50382 not n16899 ; n16899_not
g50383 not n25899 ; n25899_not
g50384 not n19797 ; n19797_not
g50385 not n18996 ; n18996_not
g50386 not n17799 ; n17799_not
g50387 not b[14] ; b[14]_not
g50388 not n15999 ; n15999_not
g50389 not n18978 ; n18978_not
g50390 not n19887 ; n19887_not
g50391 not n19878 ; n19878_not
g50392 not n18879 ; n18879_not
g50393 not n16998 ; n16998_not
g50394 not n19698 ; n19698_not
g50395 not n17889 ; n17889_not
g50396 not n19779 ; n19779_not
g50397 not n26979 ; n26979_not
g50398 not n18987 ; n18987_not
g50399 not n18888 ; n18888_not
g50400 not n26998 ; n26998_not
g50401 not b[33] ; b[33]_not
g50402 not n18979 ; n18979_not
g50403 not a[34] ; a[34]_not
g50404 not n18997 ; n18997_not
g50405 not n17998 ; n17998_not
g50406 not b[60] ; b[60]_not
g50407 not n26989 ; n26989_not
g50408 not b[51] ; b[51]_not
g50409 not n16999 ; n16999_not
g50410 not n18889 ; n18889_not
g50411 not n18898 ; n18898_not
g50412 not n19879 ; n19879_not
g50413 not n19798 ; n19798_not
g50414 not a[61] ; a[61]_not
g50415 not n25999 ; n25999_not
g50416 not n19789 ; n19789_not
g50417 not n17989 ; n17989_not
g50418 not n19897 ; n19897_not
g50419 not b[42] ; b[42]_not
g50420 not a[43] ; a[43]_not
g50421 not b[15] ; b[15]_not
g50422 not n19969 ; n19969_not
g50423 not n19978 ; n19978_not
g50424 not a[52] ; a[52]_not
g50425 not a[25] ; a[25]_not
g50426 not b[24] ; b[24]_not
g50427 not n26899 ; n26899_not
g50428 not n19699 ; n19699_not
g50429 not a[16] ; a[16]_not
g50430 not n19888 ; n19888_not
g50431 not b[25] ; b[25]_not
g50432 not n19979 ; n19979_not
g50433 not a[62] ; a[62]_not
g50434 not a[26] ; a[26]_not
g50435 not b[52] ; b[52]_not
g50436 not n18899 ; n18899_not
g50437 not n18998 ; n18998_not
g50438 not n18989 ; n18989_not
g50439 not a[17] ; a[17]_not
g50440 not n19988 ; n19988_not
g50441 not n19799 ; n19799_not
g50442 not a[44] ; a[44]_not
g50443 not b[61] ; b[61]_not
g50444 not b[16] ; b[16]_not
g50445 not a[35] ; a[35]_not
g50446 not a[53] ; a[53]_not
g50447 not n19889 ; n19889_not
g50448 not n19997 ; n19997_not
g50449 not n17999 ; n17999_not
g50450 not n26999 ; n26999_not
g50451 not b[34] ; b[34]_not
g50452 not b[43] ; b[43]_not
g50453 not b[17] ; b[17]_not
g50454 not a[54] ; a[54]_not
g50455 not b[44] ; b[44]_not
g50456 not b[62] ; b[62]_not
g50457 not b[35] ; b[35]_not
g50458 not a[18] ; a[18]_not
g50459 not a[45] ; a[45]_not
g50460 not a[36] ; a[36]_not
g50461 not b[53] ; b[53]_not
g50462 not n19998 ; n19998_not
g50463 not b[26] ; b[26]_not
g50464 not a[27] ; a[27]_not
g50465 not n18999 ; n18999_not
g50466 not n19989 ; n19989_not
g50467 not a[63] ; a[63]_not
g50468 not b[27] ; b[27]_not
g50469 not b[36] ; b[36]_not
g50470 not b[63] ; b[63]_not
g50471 not a[28] ; a[28]_not
g50472 not a[37] ; a[37]_not
g50473 not n19999 ; n19999_not
g50474 not b[45] ; b[45]_not
g50475 not a[46] ; a[46]_not
g50476 not b[54] ; b[54]_not
g50477 not a[55] ; a[55]_not
g50478 not a[19] ; a[19]_not
g50479 not b[18] ; b[18]_not
g50480 not a[38] ; a[38]_not
g50481 not a[56] ; a[56]_not
g50482 not a[47] ; a[47]_not
g50483 not b[55] ; b[55]_not
g50484 not a[29] ; a[29]_not
g50485 not b[46] ; b[46]_not
g50486 not b[28] ; b[28]_not
g50487 not b[19] ; b[19]_not
g50488 not b[37] ; b[37]_not
g50489 not b[47] ; b[47]_not
g50490 not b[29] ; b[29]_not
g50491 not b[56] ; b[56]_not
g50492 not a[48] ; a[48]_not
g50493 not a[39] ; a[39]_not
g50494 not a[57] ; a[57]_not
g50495 not b[38] ; b[38]_not
g50496 not a[58] ; a[58]_not
g50497 not a[49] ; a[49]_not
g50498 not b[39] ; b[39]_not
g50499 not b[57] ; b[57]_not
g50500 not b[48] ; b[48]_not
g50501 not a[59] ; a[59]_not
g50502 not b[58] ; b[58]_not
g50503 not b[49] ; b[49]_not
g50504 not b[59] ; b[59]_not
o f[0]
o f[1]
o f[2]
o f[3]
o f[4]
o f[5]
o f[6]
o f[7]
o f[8]
o f[9]
o f[10]
o f[11]
o f[12]
o f[13]
o f[14]
o f[15]
o f[16]
o f[17]
o f[18]
o f[19]
o f[20]
o f[21]
o f[22]
o f[23]
o f[24]
o f[25]
o f[26]
o f[27]
o f[28]
o f[29]
o f[30]
o f[31]
o f[32]
o f[33]
o f[34]
o f[35]
o f[36]
o f[37]
o f[38]
o f[39]
o f[40]
o f[41]
o f[42]
o f[43]
o f[44]
o f[45]
o f[46]
o f[47]
o f[48]
o f[49]
o f[50]
o f[51]
o f[52]
o f[53]
o f[54]
o f[55]
o f[56]
o f[57]
o f[58]
o f[59]
o f[60]
o f[61]
o f[62]
o f[63]
o f[64]
o f[65]
o f[66]
o f[67]
o f[68]
o f[69]
o f[70]
o f[71]
o f[72]
o f[73]
o f[74]
o f[75]
o f[76]
o f[77]
o f[78]
o f[79]
o f[80]
o f[81]
o f[82]
o f[83]
o f[84]
o f[85]
o f[86]
o f[87]
o f[88]
o f[89]
o f[90]
o f[91]
o f[92]
o f[93]
o f[94]
o f[95]
o f[96]
o f[97]
o f[98]
o f[99]
o f[100]
o f[101]
o f[102]
o f[103]
o f[104]
o f[105]
o f[106]
o f[107]
o f[108]
o f[109]
o f[110]
o f[111]
o f[112]
o f[113]
o f[114]
o f[115]
o f[116]
o f[117]
o f[118]
o f[119]
o f[120]
o f[121]
o f[122]
o f[123]
o f[124]
o f[125]
o f[126]
o f[127]
