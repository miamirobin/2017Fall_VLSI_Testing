name adder
i a[0]
i a[1]
i a[2]
i a[3]
i a[4]
i a[5]
i a[6]
i a[7]
i a[8]
i a[9]
i a[10]
i a[11]
i a[12]
i a[13]
i a[14]
i a[15]
i a[16]
i a[17]
i a[18]
i a[19]
i a[20]
i a[21]
i a[22]
i a[23]
i a[24]
i a[25]
i a[26]
i a[27]
i a[28]
i a[29]
i a[30]
i a[31]
i a[32]
i a[33]
i a[34]
i a[35]
i a[36]
i a[37]
i a[38]
i a[39]
i a[40]
i a[41]
i a[42]
i a[43]
i a[44]
i a[45]
i a[46]
i a[47]
i a[48]
i a[49]
i a[50]
i a[51]
i a[52]
i a[53]
i a[54]
i a[55]
i a[56]
i a[57]
i a[58]
i a[59]
i a[60]
i a[61]
i a[62]
i a[63]
i a[64]
i a[65]
i a[66]
i a[67]
i a[68]
i a[69]
i a[70]
i a[71]
i a[72]
i a[73]
i a[74]
i a[75]
i a[76]
i a[77]
i a[78]
i a[79]
i a[80]
i a[81]
i a[82]
i a[83]
i a[84]
i a[85]
i a[86]
i a[87]
i a[88]
i a[89]
i a[90]
i a[91]
i a[92]
i a[93]
i a[94]
i a[95]
i a[96]
i a[97]
i a[98]
i a[99]
i a[100]
i a[101]
i a[102]
i a[103]
i a[104]
i a[105]
i a[106]
i a[107]
i a[108]
i a[109]
i a[110]
i a[111]
i a[112]
i a[113]
i a[114]
i a[115]
i a[116]
i a[117]
i a[118]
i a[119]
i a[120]
i a[121]
i a[122]
i a[123]
i a[124]
i a[125]
i a[126]
i a[127]
i b[0]
i b[1]
i b[2]
i b[3]
i b[4]
i b[5]
i b[6]
i b[7]
i b[8]
i b[9]
i b[10]
i b[11]
i b[12]
i b[13]
i b[14]
i b[15]
i b[16]
i b[17]
i b[18]
i b[19]
i b[20]
i b[21]
i b[22]
i b[23]
i b[24]
i b[25]
i b[26]
i b[27]
i b[28]
i b[29]
i b[30]
i b[31]
i b[32]
i b[33]
i b[34]
i b[35]
i b[36]
i b[37]
i b[38]
i b[39]
i b[40]
i b[41]
i b[42]
i b[43]
i b[44]
i b[45]
i b[46]
i b[47]
i b[48]
i b[49]
i b[50]
i b[51]
i b[52]
i b[53]
i b[54]
i b[55]
i b[56]
i b[57]
i b[58]
i b[59]
i b[60]
i b[61]
i b[62]
i b[63]
i b[64]
i b[65]
i b[66]
i b[67]
i b[68]
i b[69]
i b[70]
i b[71]
i b[72]
i b[73]
i b[74]
i b[75]
i b[76]
i b[77]
i b[78]
i b[79]
i b[80]
i b[81]
i b[82]
i b[83]
i b[84]
i b[85]
i b[86]
i b[87]
i b[88]
i b[89]
i b[90]
i b[91]
i b[92]
i b[93]
i b[94]
i b[95]
i b[96]
i b[97]
i b[98]
i b[99]
i b[100]
i b[101]
i b[102]
i b[103]
i b[104]
i b[105]
i b[106]
i b[107]
i b[108]
i b[109]
i b[110]
i b[111]
i b[112]
i b[113]
i b[114]
i b[115]
i b[116]
i b[117]
i b[118]
i b[119]
i b[120]
i b[121]
i b[122]
i b[123]
i b[124]
i b[125]
i b[126]
i b[127]

g1 and a[0] b[0]_not ; n386
g2 and a[0]_not b[0] ; n387
g3 and n386_not n387_not ; f[0]
g4 and a[0] b[0] ; n389
g5 and a[1]_not b[1]_not ; n390
g6 and a[1] b[1] ; n391
g7 and n390_not n391_not ; n392
g8 and n389 n392_not ; n393
g9 and n389_not n392 ; n394
g10 and n393_not n394_not ; f[1]
g11 and n389 n390_not ; n396
g12 and n391_not n396_not ; n397
g13 and a[2]_not b[2]_not ; n398
g14 and a[2] b[2] ; n399
g15 and n398_not n399_not ; n400
g16 and n397 n400_not ; n401
g17 and n397_not n400 ; n402
g18 and n401_not n402_not ; f[2]
g19 and n397_not n398_not ; n404
g20 and n399_not n404_not ; n405
g21 and a[3]_not b[3]_not ; n406
g22 and a[3] b[3] ; n407
g23 and n406_not n407_not ; n408
g24 and n405 n408_not ; n409
g25 and n405_not n408 ; n410
g26 and n409_not n410_not ; f[3]
g27 and n405_not n406_not ; n412
g28 and n407_not n412_not ; n413
g29 and a[4]_not b[4]_not ; n414
g30 and a[4] b[4] ; n415
g31 and n414_not n415_not ; n416
g32 and n413 n416_not ; n417
g33 and n413_not n416 ; n418
g34 and n417_not n418_not ; f[4]
g35 and n413_not n414_not ; n420
g36 and n415_not n420_not ; n421
g37 and a[5]_not b[5]_not ; n422
g38 and a[5] b[5] ; n423
g39 and n422_not n423_not ; n424
g40 and n421 n424_not ; n425
g41 and n421_not n424 ; n426
g42 and n425_not n426_not ; f[5]
g43 and n421_not n422_not ; n428
g44 and n423_not n428_not ; n429
g45 and a[6]_not b[6]_not ; n430
g46 and a[6] b[6] ; n431
g47 and n430_not n431_not ; n432
g48 and n429 n432_not ; n433
g49 and n429_not n432 ; n434
g50 and n433_not n434_not ; f[6]
g51 and n429_not n430_not ; n436
g52 and n431_not n436_not ; n437
g53 and a[7]_not b[7]_not ; n438
g54 and a[7] b[7] ; n439
g55 and n438_not n439_not ; n440
g56 and n437 n440_not ; n441
g57 and n437_not n440 ; n442
g58 and n441_not n442_not ; f[7]
g59 and n437_not n438_not ; n444
g60 and n439_not n444_not ; n445
g61 and a[8]_not b[8]_not ; n446
g62 and a[8] b[8] ; n447
g63 and n446_not n447_not ; n448
g64 and n445 n448_not ; n449
g65 and n445_not n448 ; n450
g66 and n449_not n450_not ; f[8]
g67 and n445_not n446_not ; n452
g68 and n447_not n452_not ; n453
g69 and a[9]_not b[9]_not ; n454
g70 and a[9] b[9] ; n455
g71 and n454_not n455_not ; n456
g72 and n453 n456_not ; n457
g73 and n453_not n456 ; n458
g74 and n457_not n458_not ; f[9]
g75 and n453_not n454_not ; n460
g76 and n455_not n460_not ; n461
g77 and a[10]_not b[10]_not ; n462
g78 and a[10] b[10] ; n463
g79 and n462_not n463_not ; n464
g80 and n461 n464_not ; n465
g81 and n461_not n464 ; n466
g82 and n465_not n466_not ; f[10]
g83 and n461_not n462_not ; n468
g84 and n463_not n468_not ; n469
g85 and a[11]_not b[11]_not ; n470
g86 and a[11] b[11] ; n471
g87 and n470_not n471_not ; n472
g88 and n469 n472_not ; n473
g89 and n469_not n472 ; n474
g90 and n473_not n474_not ; f[11]
g91 and n469_not n470_not ; n476
g92 and n471_not n476_not ; n477
g93 and a[12]_not b[12]_not ; n478
g94 and a[12] b[12] ; n479
g95 and n478_not n479_not ; n480
g96 and n477 n480_not ; n481
g97 and n477_not n480 ; n482
g98 and n481_not n482_not ; f[12]
g99 and n477_not n478_not ; n484
g100 and n479_not n484_not ; n485
g101 and a[13]_not b[13]_not ; n486
g102 and a[13] b[13] ; n487
g103 and n486_not n487_not ; n488
g104 and n485 n488_not ; n489
g105 and n485_not n488 ; n490
g106 and n489_not n490_not ; f[13]
g107 and n485_not n486_not ; n492
g108 and n487_not n492_not ; n493
g109 and a[14]_not b[14]_not ; n494
g110 and a[14] b[14] ; n495
g111 and n494_not n495_not ; n496
g112 and n493 n496_not ; n497
g113 and n493_not n496 ; n498
g114 and n497_not n498_not ; f[14]
g115 and n493_not n494_not ; n500
g116 and n495_not n500_not ; n501
g117 and a[15]_not b[15]_not ; n502
g118 and a[15] b[15] ; n503
g119 and n502_not n503_not ; n504
g120 and n501 n504_not ; n505
g121 and n501_not n504 ; n506
g122 and n505_not n506_not ; f[15]
g123 and n501_not n502_not ; n508
g124 and n503_not n508_not ; n509
g125 and a[16]_not b[16]_not ; n510
g126 and a[16] b[16] ; n511
g127 and n510_not n511_not ; n512
g128 and n509 n512_not ; n513
g129 and n509_not n512 ; n514
g130 and n513_not n514_not ; f[16]
g131 and n509_not n510_not ; n516
g132 and n511_not n516_not ; n517
g133 and a[17]_not b[17]_not ; n518
g134 and a[17] b[17] ; n519
g135 and n518_not n519_not ; n520
g136 and n517 n520_not ; n521
g137 and n517_not n520 ; n522
g138 and n521_not n522_not ; f[17]
g139 and n517_not n518_not ; n524
g140 and n519_not n524_not ; n525
g141 and a[18]_not b[18]_not ; n526
g142 and a[18] b[18] ; n527
g143 and n526_not n527_not ; n528
g144 and n525 n528_not ; n529
g145 and n525_not n528 ; n530
g146 and n529_not n530_not ; f[18]
g147 and n525_not n526_not ; n532
g148 and n527_not n532_not ; n533
g149 and a[19]_not b[19]_not ; n534
g150 and a[19] b[19] ; n535
g151 and n534_not n535_not ; n536
g152 and n533 n536_not ; n537
g153 and n533_not n536 ; n538
g154 and n537_not n538_not ; f[19]
g155 and n533_not n534_not ; n540
g156 and n535_not n540_not ; n541
g157 and a[20]_not b[20]_not ; n542
g158 and a[20] b[20] ; n543
g159 and n542_not n543_not ; n544
g160 and n541 n544_not ; n545
g161 and n541_not n544 ; n546
g162 and n545_not n546_not ; f[20]
g163 and n541_not n542_not ; n548
g164 and n543_not n548_not ; n549
g165 and a[21]_not b[21]_not ; n550
g166 and a[21] b[21] ; n551
g167 and n550_not n551_not ; n552
g168 and n549 n552_not ; n553
g169 and n549_not n552 ; n554
g170 and n553_not n554_not ; f[21]
g171 and n549_not n550_not ; n556
g172 and n551_not n556_not ; n557
g173 and a[22]_not b[22]_not ; n558
g174 and a[22] b[22] ; n559
g175 and n558_not n559_not ; n560
g176 and n557 n560_not ; n561
g177 and n557_not n560 ; n562
g178 and n561_not n562_not ; f[22]
g179 and n557_not n558_not ; n564
g180 and n559_not n564_not ; n565
g181 and a[23]_not b[23]_not ; n566
g182 and a[23] b[23] ; n567
g183 and n566_not n567_not ; n568
g184 and n565 n568_not ; n569
g185 and n565_not n568 ; n570
g186 and n569_not n570_not ; f[23]
g187 and n565_not n566_not ; n572
g188 and n567_not n572_not ; n573
g189 and a[24]_not b[24]_not ; n574
g190 and a[24] b[24] ; n575
g191 and n574_not n575_not ; n576
g192 and n573 n576_not ; n577
g193 and n573_not n576 ; n578
g194 and n577_not n578_not ; f[24]
g195 and n573_not n574_not ; n580
g196 and n575_not n580_not ; n581
g197 and a[25]_not b[25]_not ; n582
g198 and a[25] b[25] ; n583
g199 and n582_not n583_not ; n584
g200 and n581 n584_not ; n585
g201 and n581_not n584 ; n586
g202 and n585_not n586_not ; f[25]
g203 and n581_not n582_not ; n588
g204 and n583_not n588_not ; n589
g205 and a[26]_not b[26]_not ; n590
g206 and a[26] b[26] ; n591
g207 and n590_not n591_not ; n592
g208 and n589 n592_not ; n593
g209 and n589_not n592 ; n594
g210 and n593_not n594_not ; f[26]
g211 and n589_not n590_not ; n596
g212 and n591_not n596_not ; n597
g213 and a[27]_not b[27]_not ; n598
g214 and a[27] b[27] ; n599
g215 and n598_not n599_not ; n600
g216 and n597 n600_not ; n601
g217 and n597_not n600 ; n602
g218 and n601_not n602_not ; f[27]
g219 and n597_not n598_not ; n604
g220 and n599_not n604_not ; n605
g221 and a[28]_not b[28]_not ; n606
g222 and a[28] b[28] ; n607
g223 and n606_not n607_not ; n608
g224 and n605 n608_not ; n609
g225 and n605_not n608 ; n610
g226 and n609_not n610_not ; f[28]
g227 and n605_not n606_not ; n612
g228 and n607_not n612_not ; n613
g229 and a[29]_not b[29]_not ; n614
g230 and a[29] b[29] ; n615
g231 and n614_not n615_not ; n616
g232 and n613 n616_not ; n617
g233 and n613_not n616 ; n618
g234 and n617_not n618_not ; f[29]
g235 and n613_not n614_not ; n620
g236 and n615_not n620_not ; n621
g237 and a[30]_not b[30]_not ; n622
g238 and a[30] b[30] ; n623
g239 and n622_not n623_not ; n624
g240 and n621 n624_not ; n625
g241 and n621_not n624 ; n626
g242 and n625_not n626_not ; f[30]
g243 and n621_not n622_not ; n628
g244 and n623_not n628_not ; n629
g245 and a[31]_not b[31]_not ; n630
g246 and a[31] b[31] ; n631
g247 and n630_not n631_not ; n632
g248 and n629 n632_not ; n633
g249 and n629_not n632 ; n634
g250 and n633_not n634_not ; f[31]
g251 and n629_not n630_not ; n636
g252 and n631_not n636_not ; n637
g253 and a[32]_not b[32]_not ; n638
g254 and a[32] b[32] ; n639
g255 and n638_not n639_not ; n640
g256 and n637 n640_not ; n641
g257 and n637_not n640 ; n642
g258 and n641_not n642_not ; f[32]
g259 and n637_not n638_not ; n644
g260 and n639_not n644_not ; n645
g261 and a[33]_not b[33]_not ; n646
g262 and a[33] b[33] ; n647
g263 and n646_not n647_not ; n648
g264 and n645 n648_not ; n649
g265 and n645_not n648 ; n650
g266 and n649_not n650_not ; f[33]
g267 and n645_not n646_not ; n652
g268 and n647_not n652_not ; n653
g269 and a[34]_not b[34]_not ; n654
g270 and a[34] b[34] ; n655
g271 and n654_not n655_not ; n656
g272 and n653 n656_not ; n657
g273 and n653_not n656 ; n658
g274 and n657_not n658_not ; f[34]
g275 and n653_not n654_not ; n660
g276 and n655_not n660_not ; n661
g277 and a[35]_not b[35]_not ; n662
g278 and a[35] b[35] ; n663
g279 and n662_not n663_not ; n664
g280 and n661 n664_not ; n665
g281 and n661_not n664 ; n666
g282 and n665_not n666_not ; f[35]
g283 and n661_not n662_not ; n668
g284 and n663_not n668_not ; n669
g285 and a[36]_not b[36]_not ; n670
g286 and a[36] b[36] ; n671
g287 and n670_not n671_not ; n672
g288 and n669 n672_not ; n673
g289 and n669_not n672 ; n674
g290 and n673_not n674_not ; f[36]
g291 and n669_not n670_not ; n676
g292 and n671_not n676_not ; n677
g293 and a[37]_not b[37]_not ; n678
g294 and a[37] b[37] ; n679
g295 and n678_not n679_not ; n680
g296 and n677 n680_not ; n681
g297 and n677_not n680 ; n682
g298 and n681_not n682_not ; f[37]
g299 and n677_not n678_not ; n684
g300 and n679_not n684_not ; n685
g301 and a[38]_not b[38]_not ; n686
g302 and a[38] b[38] ; n687
g303 and n686_not n687_not ; n688
g304 and n685 n688_not ; n689
g305 and n685_not n688 ; n690
g306 and n689_not n690_not ; f[38]
g307 and n685_not n686_not ; n692
g308 and n687_not n692_not ; n693
g309 and a[39]_not b[39]_not ; n694
g310 and a[39] b[39] ; n695
g311 and n694_not n695_not ; n696
g312 and n693 n696_not ; n697
g313 and n693_not n696 ; n698
g314 and n697_not n698_not ; f[39]
g315 and n693_not n694_not ; n700
g316 and n695_not n700_not ; n701
g317 and a[40]_not b[40]_not ; n702
g318 and a[40] b[40] ; n703
g319 and n702_not n703_not ; n704
g320 and n701 n704_not ; n705
g321 and n701_not n704 ; n706
g322 and n705_not n706_not ; f[40]
g323 and n701_not n702_not ; n708
g324 and n703_not n708_not ; n709
g325 and a[41]_not b[41]_not ; n710
g326 and a[41] b[41] ; n711
g327 and n710_not n711_not ; n712
g328 and n709 n712_not ; n713
g329 and n709_not n712 ; n714
g330 and n713_not n714_not ; f[41]
g331 and n709_not n710_not ; n716
g332 and n711_not n716_not ; n717
g333 and a[42]_not b[42]_not ; n718
g334 and a[42] b[42] ; n719
g335 and n718_not n719_not ; n720
g336 and n717 n720_not ; n721
g337 and n717_not n720 ; n722
g338 and n721_not n722_not ; f[42]
g339 and n717_not n718_not ; n724
g340 and n719_not n724_not ; n725
g341 and a[43]_not b[43]_not ; n726
g342 and a[43] b[43] ; n727
g343 and n726_not n727_not ; n728
g344 and n725 n728_not ; n729
g345 and n725_not n728 ; n730
g346 and n729_not n730_not ; f[43]
g347 and n725_not n726_not ; n732
g348 and n727_not n732_not ; n733
g349 and a[44]_not b[44]_not ; n734
g350 and a[44] b[44] ; n735
g351 and n734_not n735_not ; n736
g352 and n733 n736_not ; n737
g353 and n733_not n736 ; n738
g354 and n737_not n738_not ; f[44]
g355 and n733_not n734_not ; n740
g356 and n735_not n740_not ; n741
g357 and a[45]_not b[45]_not ; n742
g358 and a[45] b[45] ; n743
g359 and n742_not n743_not ; n744
g360 and n741 n744_not ; n745
g361 and n741_not n744 ; n746
g362 and n745_not n746_not ; f[45]
g363 and n741_not n742_not ; n748
g364 and n743_not n748_not ; n749
g365 and a[46]_not b[46]_not ; n750
g366 and a[46] b[46] ; n751
g367 and n750_not n751_not ; n752
g368 and n749 n752_not ; n753
g369 and n749_not n752 ; n754
g370 and n753_not n754_not ; f[46]
g371 and n749_not n750_not ; n756
g372 and n751_not n756_not ; n757
g373 and a[47]_not b[47]_not ; n758
g374 and a[47] b[47] ; n759
g375 and n758_not n759_not ; n760
g376 and n757 n760_not ; n761
g377 and n757_not n760 ; n762
g378 and n761_not n762_not ; f[47]
g379 and n757_not n758_not ; n764
g380 and n759_not n764_not ; n765
g381 and a[48]_not b[48]_not ; n766
g382 and a[48] b[48] ; n767
g383 and n766_not n767_not ; n768
g384 and n765 n768_not ; n769
g385 and n765_not n768 ; n770
g386 and n769_not n770_not ; f[48]
g387 and n765_not n766_not ; n772
g388 and n767_not n772_not ; n773
g389 and a[49]_not b[49]_not ; n774
g390 and a[49] b[49] ; n775
g391 and n774_not n775_not ; n776
g392 and n773 n776_not ; n777
g393 and n773_not n776 ; n778
g394 and n777_not n778_not ; f[49]
g395 and n773_not n774_not ; n780
g396 and n775_not n780_not ; n781
g397 and a[50]_not b[50]_not ; n782
g398 and a[50] b[50] ; n783
g399 and n782_not n783_not ; n784
g400 and n781 n784_not ; n785
g401 and n781_not n784 ; n786
g402 and n785_not n786_not ; f[50]
g403 and n781_not n782_not ; n788
g404 and n783_not n788_not ; n789
g405 and a[51]_not b[51]_not ; n790
g406 and a[51] b[51] ; n791
g407 and n790_not n791_not ; n792
g408 and n789 n792_not ; n793
g409 and n789_not n792 ; n794
g410 and n793_not n794_not ; f[51]
g411 and n789_not n790_not ; n796
g412 and n791_not n796_not ; n797
g413 and a[52]_not b[52]_not ; n798
g414 and a[52] b[52] ; n799
g415 and n798_not n799_not ; n800
g416 and n797 n800_not ; n801
g417 and n797_not n800 ; n802
g418 and n801_not n802_not ; f[52]
g419 and n797_not n798_not ; n804
g420 and n799_not n804_not ; n805
g421 and a[53]_not b[53]_not ; n806
g422 and a[53] b[53] ; n807
g423 and n806_not n807_not ; n808
g424 and n805 n808_not ; n809
g425 and n805_not n808 ; n810
g426 and n809_not n810_not ; f[53]
g427 and n805_not n806_not ; n812
g428 and n807_not n812_not ; n813
g429 and a[54]_not b[54]_not ; n814
g430 and a[54] b[54] ; n815
g431 and n814_not n815_not ; n816
g432 and n813 n816_not ; n817
g433 and n813_not n816 ; n818
g434 and n817_not n818_not ; f[54]
g435 and n813_not n814_not ; n820
g436 and n815_not n820_not ; n821
g437 and a[55]_not b[55]_not ; n822
g438 and a[55] b[55] ; n823
g439 and n822_not n823_not ; n824
g440 and n821 n824_not ; n825
g441 and n821_not n824 ; n826
g442 and n825_not n826_not ; f[55]
g443 and n821_not n822_not ; n828
g444 and n823_not n828_not ; n829
g445 and a[56]_not b[56]_not ; n830
g446 and a[56] b[56] ; n831
g447 and n830_not n831_not ; n832
g448 and n829 n832_not ; n833
g449 and n829_not n832 ; n834
g450 and n833_not n834_not ; f[56]
g451 and n829_not n830_not ; n836
g452 and n831_not n836_not ; n837
g453 and a[57]_not b[57]_not ; n838
g454 and a[57] b[57] ; n839
g455 and n838_not n839_not ; n840
g456 and n837 n840_not ; n841
g457 and n837_not n840 ; n842
g458 and n841_not n842_not ; f[57]
g459 and n837_not n838_not ; n844
g460 and n839_not n844_not ; n845
g461 and a[58]_not b[58]_not ; n846
g462 and a[58] b[58] ; n847
g463 and n846_not n847_not ; n848
g464 and n845 n848_not ; n849
g465 and n845_not n848 ; n850
g466 and n849_not n850_not ; f[58]
g467 and n845_not n846_not ; n852
g468 and n847_not n852_not ; n853
g469 and a[59]_not b[59]_not ; n854
g470 and a[59] b[59] ; n855
g471 and n854_not n855_not ; n856
g472 and n853 n856_not ; n857
g473 and n853_not n856 ; n858
g474 and n857_not n858_not ; f[59]
g475 and n853_not n854_not ; n860
g476 and n855_not n860_not ; n861
g477 and a[60]_not b[60]_not ; n862
g478 and a[60] b[60] ; n863
g479 and n862_not n863_not ; n864
g480 and n861 n864_not ; n865
g481 and n861_not n864 ; n866
g482 and n865_not n866_not ; f[60]
g483 and n861_not n862_not ; n868
g484 and n863_not n868_not ; n869
g485 and a[61]_not b[61]_not ; n870
g486 and a[61] b[61] ; n871
g487 and n870_not n871_not ; n872
g488 and n869 n872_not ; n873
g489 and n869_not n872 ; n874
g490 and n873_not n874_not ; f[61]
g491 and n869_not n870_not ; n876
g492 and n871_not n876_not ; n877
g493 and a[62]_not b[62]_not ; n878
g494 and a[62] b[62] ; n879
g495 and n878_not n879_not ; n880
g496 and n877 n880_not ; n881
g497 and n877_not n880 ; n882
g498 and n881_not n882_not ; f[62]
g499 and n877_not n878_not ; n884
g500 and n879_not n884_not ; n885
g501 and a[63]_not b[63]_not ; n886
g502 and a[63] b[63] ; n887
g503 and n886_not n887_not ; n888
g504 and n885 n888_not ; n889
g505 and n885_not n888 ; n890
g506 and n889_not n890_not ; f[63]
g507 and n885_not n886_not ; n892
g508 and n887_not n892_not ; n893
g509 and a[64]_not b[64]_not ; n894
g510 and a[64] b[64] ; n895
g511 and n894_not n895_not ; n896
g512 and n893 n896_not ; n897
g513 and n893_not n896 ; n898
g514 and n897_not n898_not ; f[64]
g515 and n893_not n894_not ; n900
g516 and n895_not n900_not ; n901
g517 and a[65]_not b[65]_not ; n902
g518 and a[65] b[65] ; n903
g519 and n902_not n903_not ; n904
g520 and n901 n904_not ; n905
g521 and n901_not n904 ; n906
g522 and n905_not n906_not ; f[65]
g523 and n901_not n902_not ; n908
g524 and n903_not n908_not ; n909
g525 and a[66]_not b[66]_not ; n910
g526 and a[66] b[66] ; n911
g527 and n910_not n911_not ; n912
g528 and n909 n912_not ; n913
g529 and n909_not n912 ; n914
g530 and n913_not n914_not ; f[66]
g531 and n909_not n910_not ; n916
g532 and n911_not n916_not ; n917
g533 and a[67]_not b[67]_not ; n918
g534 and a[67] b[67] ; n919
g535 and n918_not n919_not ; n920
g536 and n917 n920_not ; n921
g537 and n917_not n920 ; n922
g538 and n921_not n922_not ; f[67]
g539 and n917_not n918_not ; n924
g540 and n919_not n924_not ; n925
g541 and a[68]_not b[68]_not ; n926
g542 and a[68] b[68] ; n927
g543 and n926_not n927_not ; n928
g544 and n925 n928_not ; n929
g545 and n925_not n928 ; n930
g546 and n929_not n930_not ; f[68]
g547 and n925_not n926_not ; n932
g548 and n927_not n932_not ; n933
g549 and a[69]_not b[69]_not ; n934
g550 and a[69] b[69] ; n935
g551 and n934_not n935_not ; n936
g552 and n933 n936_not ; n937
g553 and n933_not n936 ; n938
g554 and n937_not n938_not ; f[69]
g555 and n933_not n934_not ; n940
g556 and n935_not n940_not ; n941
g557 and a[70]_not b[70]_not ; n942
g558 and a[70] b[70] ; n943
g559 and n942_not n943_not ; n944
g560 and n941 n944_not ; n945
g561 and n941_not n944 ; n946
g562 and n945_not n946_not ; f[70]
g563 and n941_not n942_not ; n948
g564 and n943_not n948_not ; n949
g565 and a[71]_not b[71]_not ; n950
g566 and a[71] b[71] ; n951
g567 and n950_not n951_not ; n952
g568 and n949 n952_not ; n953
g569 and n949_not n952 ; n954
g570 and n953_not n954_not ; f[71]
g571 and n949_not n950_not ; n956
g572 and n951_not n956_not ; n957
g573 and a[72]_not b[72]_not ; n958
g574 and a[72] b[72] ; n959
g575 and n958_not n959_not ; n960
g576 and n957 n960_not ; n961
g577 and n957_not n960 ; n962
g578 and n961_not n962_not ; f[72]
g579 and n957_not n958_not ; n964
g580 and n959_not n964_not ; n965
g581 and a[73]_not b[73]_not ; n966
g582 and a[73] b[73] ; n967
g583 and n966_not n967_not ; n968
g584 and n965 n968_not ; n969
g585 and n965_not n968 ; n970
g586 and n969_not n970_not ; f[73]
g587 and n965_not n966_not ; n972
g588 and n967_not n972_not ; n973
g589 and a[74]_not b[74]_not ; n974
g590 and a[74] b[74] ; n975
g591 and n974_not n975_not ; n976
g592 and n973 n976_not ; n977
g593 and n973_not n976 ; n978
g594 and n977_not n978_not ; f[74]
g595 and n973_not n974_not ; n980
g596 and n975_not n980_not ; n981
g597 and a[75]_not b[75]_not ; n982
g598 and a[75] b[75] ; n983
g599 and n982_not n983_not ; n984
g600 and n981 n984_not ; n985
g601 and n981_not n984 ; n986
g602 and n985_not n986_not ; f[75]
g603 and n981_not n982_not ; n988
g604 and n983_not n988_not ; n989
g605 and a[76]_not b[76]_not ; n990
g606 and a[76] b[76] ; n991
g607 and n990_not n991_not ; n992
g608 and n989 n992_not ; n993
g609 and n989_not n992 ; n994
g610 and n993_not n994_not ; f[76]
g611 and n989_not n990_not ; n996
g612 and n991_not n996_not ; n997
g613 and a[77]_not b[77]_not ; n998
g614 and a[77] b[77] ; n999
g615 and n998_not n999_not ; n1000
g616 and n997 n1000_not ; n1001
g617 and n997_not n1000 ; n1002
g618 and n1001_not n1002_not ; f[77]
g619 and n997_not n998_not ; n1004
g620 and n999_not n1004_not ; n1005
g621 and a[78]_not b[78]_not ; n1006
g622 and a[78] b[78] ; n1007
g623 and n1006_not n1007_not ; n1008
g624 and n1005 n1008_not ; n1009
g625 and n1005_not n1008 ; n1010
g626 and n1009_not n1010_not ; f[78]
g627 and n1005_not n1006_not ; n1012
g628 and n1007_not n1012_not ; n1013
g629 and a[79]_not b[79]_not ; n1014
g630 and a[79] b[79] ; n1015
g631 and n1014_not n1015_not ; n1016
g632 and n1013 n1016_not ; n1017
g633 and n1013_not n1016 ; n1018
g634 and n1017_not n1018_not ; f[79]
g635 and n1013_not n1014_not ; n1020
g636 and n1015_not n1020_not ; n1021
g637 and a[80]_not b[80]_not ; n1022
g638 and a[80] b[80] ; n1023
g639 and n1022_not n1023_not ; n1024
g640 and n1021 n1024_not ; n1025
g641 and n1021_not n1024 ; n1026
g642 and n1025_not n1026_not ; f[80]
g643 and n1021_not n1022_not ; n1028
g644 and n1023_not n1028_not ; n1029
g645 and a[81]_not b[81]_not ; n1030
g646 and a[81] b[81] ; n1031
g647 and n1030_not n1031_not ; n1032
g648 and n1029 n1032_not ; n1033
g649 and n1029_not n1032 ; n1034
g650 and n1033_not n1034_not ; f[81]
g651 and n1029_not n1030_not ; n1036
g652 and n1031_not n1036_not ; n1037
g653 and a[82]_not b[82]_not ; n1038
g654 and a[82] b[82] ; n1039
g655 and n1038_not n1039_not ; n1040
g656 and n1037 n1040_not ; n1041
g657 and n1037_not n1040 ; n1042
g658 and n1041_not n1042_not ; f[82]
g659 and n1037_not n1038_not ; n1044
g660 and n1039_not n1044_not ; n1045
g661 and a[83]_not b[83]_not ; n1046
g662 and a[83] b[83] ; n1047
g663 and n1046_not n1047_not ; n1048
g664 and n1045 n1048_not ; n1049
g665 and n1045_not n1048 ; n1050
g666 and n1049_not n1050_not ; f[83]
g667 and n1045_not n1046_not ; n1052
g668 and n1047_not n1052_not ; n1053
g669 and a[84]_not b[84]_not ; n1054
g670 and a[84] b[84] ; n1055
g671 and n1054_not n1055_not ; n1056
g672 and n1053 n1056_not ; n1057
g673 and n1053_not n1056 ; n1058
g674 and n1057_not n1058_not ; f[84]
g675 and n1053_not n1054_not ; n1060
g676 and n1055_not n1060_not ; n1061
g677 and a[85]_not b[85]_not ; n1062
g678 and a[85] b[85] ; n1063
g679 and n1062_not n1063_not ; n1064
g680 and n1061 n1064_not ; n1065
g681 and n1061_not n1064 ; n1066
g682 and n1065_not n1066_not ; f[85]
g683 and n1061_not n1062_not ; n1068
g684 and n1063_not n1068_not ; n1069
g685 and a[86]_not b[86]_not ; n1070
g686 and a[86] b[86] ; n1071
g687 and n1070_not n1071_not ; n1072
g688 and n1069 n1072_not ; n1073
g689 and n1069_not n1072 ; n1074
g690 and n1073_not n1074_not ; f[86]
g691 and n1069_not n1070_not ; n1076
g692 and n1071_not n1076_not ; n1077
g693 and a[87]_not b[87]_not ; n1078
g694 and a[87] b[87] ; n1079
g695 and n1078_not n1079_not ; n1080
g696 and n1077 n1080_not ; n1081
g697 and n1077_not n1080 ; n1082
g698 and n1081_not n1082_not ; f[87]
g699 and n1077_not n1078_not ; n1084
g700 and n1079_not n1084_not ; n1085
g701 and a[88]_not b[88]_not ; n1086
g702 and a[88] b[88] ; n1087
g703 and n1086_not n1087_not ; n1088
g704 and n1085 n1088_not ; n1089
g705 and n1085_not n1088 ; n1090
g706 and n1089_not n1090_not ; f[88]
g707 and n1085_not n1086_not ; n1092
g708 and n1087_not n1092_not ; n1093
g709 and a[89]_not b[89]_not ; n1094
g710 and a[89] b[89] ; n1095
g711 and n1094_not n1095_not ; n1096
g712 and n1093 n1096_not ; n1097
g713 and n1093_not n1096 ; n1098
g714 and n1097_not n1098_not ; f[89]
g715 and n1093_not n1094_not ; n1100
g716 and n1095_not n1100_not ; n1101
g717 and a[90]_not b[90]_not ; n1102
g718 and a[90] b[90] ; n1103
g719 and n1102_not n1103_not ; n1104
g720 and n1101 n1104_not ; n1105
g721 and n1101_not n1104 ; n1106
g722 and n1105_not n1106_not ; f[90]
g723 and n1101_not n1102_not ; n1108
g724 and n1103_not n1108_not ; n1109
g725 and a[91]_not b[91]_not ; n1110
g726 and a[91] b[91] ; n1111
g727 and n1110_not n1111_not ; n1112
g728 and n1109 n1112_not ; n1113
g729 and n1109_not n1112 ; n1114
g730 and n1113_not n1114_not ; f[91]
g731 and n1109_not n1110_not ; n1116
g732 and n1111_not n1116_not ; n1117
g733 and a[92]_not b[92]_not ; n1118
g734 and a[92] b[92] ; n1119
g735 and n1118_not n1119_not ; n1120
g736 and n1117 n1120_not ; n1121
g737 and n1117_not n1120 ; n1122
g738 and n1121_not n1122_not ; f[92]
g739 and n1117_not n1118_not ; n1124
g740 and n1119_not n1124_not ; n1125
g741 and a[93]_not b[93]_not ; n1126
g742 and a[93] b[93] ; n1127
g743 and n1126_not n1127_not ; n1128
g744 and n1125 n1128_not ; n1129
g745 and n1125_not n1128 ; n1130
g746 and n1129_not n1130_not ; f[93]
g747 and n1125_not n1126_not ; n1132
g748 and n1127_not n1132_not ; n1133
g749 and a[94]_not b[94]_not ; n1134
g750 and a[94] b[94] ; n1135
g751 and n1134_not n1135_not ; n1136
g752 and n1133 n1136_not ; n1137
g753 and n1133_not n1136 ; n1138
g754 and n1137_not n1138_not ; f[94]
g755 and n1133_not n1134_not ; n1140
g756 and n1135_not n1140_not ; n1141
g757 and a[95]_not b[95]_not ; n1142
g758 and a[95] b[95] ; n1143
g759 and n1142_not n1143_not ; n1144
g760 and n1141 n1144_not ; n1145
g761 and n1141_not n1144 ; n1146
g762 and n1145_not n1146_not ; f[95]
g763 and n1141_not n1142_not ; n1148
g764 and n1143_not n1148_not ; n1149
g765 and a[96]_not b[96]_not ; n1150
g766 and a[96] b[96] ; n1151
g767 and n1150_not n1151_not ; n1152
g768 and n1149 n1152_not ; n1153
g769 and n1149_not n1152 ; n1154
g770 and n1153_not n1154_not ; f[96]
g771 and n1149_not n1150_not ; n1156
g772 and n1151_not n1156_not ; n1157
g773 and a[97]_not b[97]_not ; n1158
g774 and a[97] b[97] ; n1159
g775 and n1158_not n1159_not ; n1160
g776 and n1157 n1160_not ; n1161
g777 and n1157_not n1160 ; n1162
g778 and n1161_not n1162_not ; f[97]
g779 and n1157_not n1158_not ; n1164
g780 and n1159_not n1164_not ; n1165
g781 and a[98]_not b[98]_not ; n1166
g782 and a[98] b[98] ; n1167
g783 and n1166_not n1167_not ; n1168
g784 and n1165 n1168_not ; n1169
g785 and n1165_not n1168 ; n1170
g786 and n1169_not n1170_not ; f[98]
g787 and n1165_not n1166_not ; n1172
g788 and n1167_not n1172_not ; n1173
g789 and a[99]_not b[99]_not ; n1174
g790 and a[99] b[99] ; n1175
g791 and n1174_not n1175_not ; n1176
g792 and n1173 n1176_not ; n1177
g793 and n1173_not n1176 ; n1178
g794 and n1177_not n1178_not ; f[99]
g795 and n1173_not n1174_not ; n1180
g796 and n1175_not n1180_not ; n1181
g797 and a[100]_not b[100]_not ; n1182
g798 and a[100] b[100] ; n1183
g799 and n1182_not n1183_not ; n1184
g800 and n1181 n1184_not ; n1185
g801 and n1181_not n1184 ; n1186
g802 and n1185_not n1186_not ; f[100]
g803 and n1181_not n1182_not ; n1188
g804 and n1183_not n1188_not ; n1189
g805 and a[101]_not b[101]_not ; n1190
g806 and a[101] b[101] ; n1191
g807 and n1190_not n1191_not ; n1192
g808 and n1189 n1192_not ; n1193
g809 and n1189_not n1192 ; n1194
g810 and n1193_not n1194_not ; f[101]
g811 and n1189_not n1190_not ; n1196
g812 and n1191_not n1196_not ; n1197
g813 and a[102]_not b[102]_not ; n1198
g814 and a[102] b[102] ; n1199
g815 and n1198_not n1199_not ; n1200
g816 and n1197 n1200_not ; n1201
g817 and n1197_not n1200 ; n1202
g818 and n1201_not n1202_not ; f[102]
g819 and n1197_not n1198_not ; n1204
g820 and n1199_not n1204_not ; n1205
g821 and a[103]_not b[103]_not ; n1206
g822 and a[103] b[103] ; n1207
g823 and n1206_not n1207_not ; n1208
g824 and n1205 n1208_not ; n1209
g825 and n1205_not n1208 ; n1210
g826 and n1209_not n1210_not ; f[103]
g827 and n1205_not n1206_not ; n1212
g828 and n1207_not n1212_not ; n1213
g829 and a[104]_not b[104]_not ; n1214
g830 and a[104] b[104] ; n1215
g831 and n1214_not n1215_not ; n1216
g832 and n1213 n1216_not ; n1217
g833 and n1213_not n1216 ; n1218
g834 and n1217_not n1218_not ; f[104]
g835 and n1213_not n1214_not ; n1220
g836 and n1215_not n1220_not ; n1221
g837 and a[105]_not b[105]_not ; n1222
g838 and a[105] b[105] ; n1223
g839 and n1222_not n1223_not ; n1224
g840 and n1221 n1224_not ; n1225
g841 and n1221_not n1224 ; n1226
g842 and n1225_not n1226_not ; f[105]
g843 and n1221_not n1222_not ; n1228
g844 and n1223_not n1228_not ; n1229
g845 and a[106]_not b[106]_not ; n1230
g846 and a[106] b[106] ; n1231
g847 and n1230_not n1231_not ; n1232
g848 and n1229 n1232_not ; n1233
g849 and n1229_not n1232 ; n1234
g850 and n1233_not n1234_not ; f[106]
g851 and n1229_not n1230_not ; n1236
g852 and n1231_not n1236_not ; n1237
g853 and a[107]_not b[107]_not ; n1238
g854 and a[107] b[107] ; n1239
g855 and n1238_not n1239_not ; n1240
g856 and n1237 n1240_not ; n1241
g857 and n1237_not n1240 ; n1242
g858 and n1241_not n1242_not ; f[107]
g859 and n1237_not n1238_not ; n1244
g860 and n1239_not n1244_not ; n1245
g861 and a[108]_not b[108]_not ; n1246
g862 and a[108] b[108] ; n1247
g863 and n1246_not n1247_not ; n1248
g864 and n1245 n1248_not ; n1249
g865 and n1245_not n1248 ; n1250
g866 and n1249_not n1250_not ; f[108]
g867 and n1245_not n1246_not ; n1252
g868 and n1247_not n1252_not ; n1253
g869 and a[109]_not b[109]_not ; n1254
g870 and a[109] b[109] ; n1255
g871 and n1254_not n1255_not ; n1256
g872 and n1253 n1256_not ; n1257
g873 and n1253_not n1256 ; n1258
g874 and n1257_not n1258_not ; f[109]
g875 and n1253_not n1254_not ; n1260
g876 and n1255_not n1260_not ; n1261
g877 and a[110]_not b[110]_not ; n1262
g878 and a[110] b[110] ; n1263
g879 and n1262_not n1263_not ; n1264
g880 and n1261 n1264_not ; n1265
g881 and n1261_not n1264 ; n1266
g882 and n1265_not n1266_not ; f[110]
g883 and n1261_not n1262_not ; n1268
g884 and n1263_not n1268_not ; n1269
g885 and a[111]_not b[111]_not ; n1270
g886 and a[111] b[111] ; n1271
g887 and n1270_not n1271_not ; n1272
g888 and n1269 n1272_not ; n1273
g889 and n1269_not n1272 ; n1274
g890 and n1273_not n1274_not ; f[111]
g891 and n1269_not n1270_not ; n1276
g892 and n1271_not n1276_not ; n1277
g893 and a[112]_not b[112]_not ; n1278
g894 and a[112] b[112] ; n1279
g895 and n1278_not n1279_not ; n1280
g896 and n1277 n1280_not ; n1281
g897 and n1277_not n1280 ; n1282
g898 and n1281_not n1282_not ; f[112]
g899 and n1277_not n1278_not ; n1284
g900 and n1279_not n1284_not ; n1285
g901 and a[113]_not b[113]_not ; n1286
g902 and a[113] b[113] ; n1287
g903 and n1286_not n1287_not ; n1288
g904 and n1285 n1288_not ; n1289
g905 and n1285_not n1288 ; n1290
g906 and n1289_not n1290_not ; f[113]
g907 and n1285_not n1286_not ; n1292
g908 and n1287_not n1292_not ; n1293
g909 and a[114]_not b[114]_not ; n1294
g910 and a[114] b[114] ; n1295
g911 and n1294_not n1295_not ; n1296
g912 and n1293 n1296_not ; n1297
g913 and n1293_not n1296 ; n1298
g914 and n1297_not n1298_not ; f[114]
g915 and n1293_not n1294_not ; n1300
g916 and n1295_not n1300_not ; n1301
g917 and a[115]_not b[115]_not ; n1302
g918 and a[115] b[115] ; n1303
g919 and n1302_not n1303_not ; n1304
g920 and n1301 n1304_not ; n1305
g921 and n1301_not n1304 ; n1306
g922 and n1305_not n1306_not ; f[115]
g923 and n1301_not n1302_not ; n1308
g924 and n1303_not n1308_not ; n1309
g925 and a[116]_not b[116]_not ; n1310
g926 and a[116] b[116] ; n1311
g927 and n1310_not n1311_not ; n1312
g928 and n1309 n1312_not ; n1313
g929 and n1309_not n1312 ; n1314
g930 and n1313_not n1314_not ; f[116]
g931 and n1309_not n1310_not ; n1316
g932 and n1311_not n1316_not ; n1317
g933 and a[117]_not b[117]_not ; n1318
g934 and a[117] b[117] ; n1319
g935 and n1318_not n1319_not ; n1320
g936 and n1317 n1320_not ; n1321
g937 and n1317_not n1320 ; n1322
g938 and n1321_not n1322_not ; f[117]
g939 and n1317_not n1318_not ; n1324
g940 and n1319_not n1324_not ; n1325
g941 and a[118]_not b[118]_not ; n1326
g942 and a[118] b[118] ; n1327
g943 and n1326_not n1327_not ; n1328
g944 and n1325 n1328_not ; n1329
g945 and n1325_not n1328 ; n1330
g946 and n1329_not n1330_not ; f[118]
g947 and n1325_not n1326_not ; n1332
g948 and n1327_not n1332_not ; n1333
g949 and a[119]_not b[119]_not ; n1334
g950 and a[119] b[119] ; n1335
g951 and n1334_not n1335_not ; n1336
g952 and n1333 n1336_not ; n1337
g953 and n1333_not n1336 ; n1338
g954 and n1337_not n1338_not ; f[119]
g955 and n1333_not n1334_not ; n1340
g956 and n1335_not n1340_not ; n1341
g957 and a[120]_not b[120]_not ; n1342
g958 and a[120] b[120] ; n1343
g959 and n1342_not n1343_not ; n1344
g960 and n1341 n1344_not ; n1345
g961 and n1341_not n1344 ; n1346
g962 and n1345_not n1346_not ; f[120]
g963 and n1341_not n1342_not ; n1348
g964 and n1343_not n1348_not ; n1349
g965 and a[121]_not b[121]_not ; n1350
g966 and a[121] b[121] ; n1351
g967 and n1350_not n1351_not ; n1352
g968 and n1349 n1352_not ; n1353
g969 and n1349_not n1352 ; n1354
g970 and n1353_not n1354_not ; f[121]
g971 and n1349_not n1350_not ; n1356
g972 and n1351_not n1356_not ; n1357
g973 and a[122]_not b[122]_not ; n1358
g974 and a[122] b[122] ; n1359
g975 and n1358_not n1359_not ; n1360
g976 and n1357 n1360_not ; n1361
g977 and n1357_not n1360 ; n1362
g978 and n1361_not n1362_not ; f[122]
g979 and n1357_not n1358_not ; n1364
g980 and n1359_not n1364_not ; n1365
g981 and a[123]_not b[123]_not ; n1366
g982 and a[123] b[123] ; n1367
g983 and n1366_not n1367_not ; n1368
g984 and n1365 n1368_not ; n1369
g985 and n1365_not n1368 ; n1370
g986 and n1369_not n1370_not ; f[123]
g987 and n1365_not n1366_not ; n1372
g988 and n1367_not n1372_not ; n1373
g989 and a[124]_not b[124]_not ; n1374
g990 and a[124] b[124] ; n1375
g991 and n1374_not n1375_not ; n1376
g992 and n1373 n1376_not ; n1377
g993 and n1373_not n1376 ; n1378
g994 and n1377_not n1378_not ; f[124]
g995 and n1373_not n1374_not ; n1380
g996 and n1375_not n1380_not ; n1381
g997 and a[125]_not b[125]_not ; n1382
g998 and a[125] b[125] ; n1383
g999 and n1382_not n1383_not ; n1384
g1000 and n1381 n1384_not ; n1385
g1001 and n1381_not n1384 ; n1386
g1002 and n1385_not n1386_not ; f[125]
g1003 and n1381_not n1382_not ; n1388
g1004 and n1383_not n1388_not ; n1389
g1005 and a[126]_not b[126]_not ; n1390
g1006 and a[126] b[126] ; n1391
g1007 and n1390_not n1391_not ; n1392
g1008 and n1389 n1392_not ; n1393
g1009 and n1389_not n1392 ; n1394
g1010 and n1393_not n1394_not ; f[126]
g1011 and n1389_not n1390_not ; n1396
g1012 and n1391_not n1396_not ; n1397
g1013 and a[127]_not b[127]_not ; n1398
g1014 and a[127] b[127] ; n1399
g1015 and n1398_not n1399_not ; n1400
g1016 and n1397 n1400_not ; n1401
g1017 and n1397_not n1400 ; n1402
g1018 and n1401_not n1402_not ; f[127]
g1019 and n1397_not n1398_not ; n1404
g1020 and n1399_not n1404_not ; cOut
g1021 not b[0] ; b[0]_not
g1022 not a[0] ; a[0]_not
g1023 not n386 ; n386_not
g1024 not n387 ; n387_not
g1025 not a[1] ; a[1]_not
g1026 not b[1] ; b[1]_not
g1027 not n390 ; n390_not
g1028 not n391 ; n391_not
g1029 not n392 ; n392_not
g1030 not n389 ; n389_not
g1031 not n393 ; n393_not
g1032 not n394 ; n394_not
g1033 not n396 ; n396_not
g1034 not a[2] ; a[2]_not
g1035 not b[2] ; b[2]_not
g1036 not n398 ; n398_not
g1037 not n399 ; n399_not
g1038 not n400 ; n400_not
g1039 not n397 ; n397_not
g1040 not n401 ; n401_not
g1041 not n402 ; n402_not
g1042 not n404 ; n404_not
g1043 not a[3] ; a[3]_not
g1044 not b[3] ; b[3]_not
g1045 not n406 ; n406_not
g1046 not n407 ; n407_not
g1047 not n408 ; n408_not
g1048 not n405 ; n405_not
g1049 not n409 ; n409_not
g1050 not n410 ; n410_not
g1051 not n412 ; n412_not
g1052 not a[4] ; a[4]_not
g1053 not b[4] ; b[4]_not
g1054 not n414 ; n414_not
g1055 not n415 ; n415_not
g1056 not n416 ; n416_not
g1057 not n413 ; n413_not
g1058 not n417 ; n417_not
g1059 not n418 ; n418_not
g1060 not n420 ; n420_not
g1061 not a[5] ; a[5]_not
g1062 not b[5] ; b[5]_not
g1063 not n422 ; n422_not
g1064 not n423 ; n423_not
g1065 not n424 ; n424_not
g1066 not n421 ; n421_not
g1067 not n425 ; n425_not
g1068 not n426 ; n426_not
g1069 not n428 ; n428_not
g1070 not a[6] ; a[6]_not
g1071 not b[6] ; b[6]_not
g1072 not n430 ; n430_not
g1073 not n431 ; n431_not
g1074 not n432 ; n432_not
g1075 not n429 ; n429_not
g1076 not n433 ; n433_not
g1077 not n434 ; n434_not
g1078 not n436 ; n436_not
g1079 not a[7] ; a[7]_not
g1080 not b[7] ; b[7]_not
g1081 not n438 ; n438_not
g1082 not n439 ; n439_not
g1083 not n440 ; n440_not
g1084 not n437 ; n437_not
g1085 not n441 ; n441_not
g1086 not n442 ; n442_not
g1087 not n444 ; n444_not
g1088 not a[8] ; a[8]_not
g1089 not b[8] ; b[8]_not
g1090 not n446 ; n446_not
g1091 not n447 ; n447_not
g1092 not n448 ; n448_not
g1093 not n445 ; n445_not
g1094 not n449 ; n449_not
g1095 not n450 ; n450_not
g1096 not n452 ; n452_not
g1097 not a[9] ; a[9]_not
g1098 not b[9] ; b[9]_not
g1099 not n454 ; n454_not
g1100 not n455 ; n455_not
g1101 not n456 ; n456_not
g1102 not n453 ; n453_not
g1103 not n457 ; n457_not
g1104 not n458 ; n458_not
g1105 not n460 ; n460_not
g1106 not a[10] ; a[10]_not
g1107 not b[10] ; b[10]_not
g1108 not n462 ; n462_not
g1109 not n463 ; n463_not
g1110 not n464 ; n464_not
g1111 not n461 ; n461_not
g1112 not n465 ; n465_not
g1113 not n466 ; n466_not
g1114 not n468 ; n468_not
g1115 not a[11] ; a[11]_not
g1116 not b[11] ; b[11]_not
g1117 not n470 ; n470_not
g1118 not n471 ; n471_not
g1119 not n472 ; n472_not
g1120 not n469 ; n469_not
g1121 not n473 ; n473_not
g1122 not n474 ; n474_not
g1123 not n476 ; n476_not
g1124 not a[12] ; a[12]_not
g1125 not b[12] ; b[12]_not
g1126 not n478 ; n478_not
g1127 not n479 ; n479_not
g1128 not n480 ; n480_not
g1129 not n477 ; n477_not
g1130 not n481 ; n481_not
g1131 not n482 ; n482_not
g1132 not n484 ; n484_not
g1133 not a[13] ; a[13]_not
g1134 not b[13] ; b[13]_not
g1135 not n486 ; n486_not
g1136 not n487 ; n487_not
g1137 not n488 ; n488_not
g1138 not n485 ; n485_not
g1139 not n489 ; n489_not
g1140 not n490 ; n490_not
g1141 not n492 ; n492_not
g1142 not a[14] ; a[14]_not
g1143 not b[14] ; b[14]_not
g1144 not n494 ; n494_not
g1145 not n495 ; n495_not
g1146 not n496 ; n496_not
g1147 not n493 ; n493_not
g1148 not n497 ; n497_not
g1149 not n498 ; n498_not
g1150 not n500 ; n500_not
g1151 not a[15] ; a[15]_not
g1152 not b[15] ; b[15]_not
g1153 not n502 ; n502_not
g1154 not n503 ; n503_not
g1155 not n504 ; n504_not
g1156 not n501 ; n501_not
g1157 not n505 ; n505_not
g1158 not n506 ; n506_not
g1159 not n508 ; n508_not
g1160 not a[16] ; a[16]_not
g1161 not b[16] ; b[16]_not
g1162 not n510 ; n510_not
g1163 not n511 ; n511_not
g1164 not n512 ; n512_not
g1165 not n509 ; n509_not
g1166 not n513 ; n513_not
g1167 not n514 ; n514_not
g1168 not n516 ; n516_not
g1169 not a[17] ; a[17]_not
g1170 not b[17] ; b[17]_not
g1171 not n518 ; n518_not
g1172 not n519 ; n519_not
g1173 not n520 ; n520_not
g1174 not n517 ; n517_not
g1175 not n521 ; n521_not
g1176 not n522 ; n522_not
g1177 not n524 ; n524_not
g1178 not a[18] ; a[18]_not
g1179 not b[18] ; b[18]_not
g1180 not n526 ; n526_not
g1181 not n527 ; n527_not
g1182 not n528 ; n528_not
g1183 not n525 ; n525_not
g1184 not n529 ; n529_not
g1185 not n530 ; n530_not
g1186 not n532 ; n532_not
g1187 not a[19] ; a[19]_not
g1188 not b[19] ; b[19]_not
g1189 not n534 ; n534_not
g1190 not n535 ; n535_not
g1191 not n536 ; n536_not
g1192 not n533 ; n533_not
g1193 not n537 ; n537_not
g1194 not n538 ; n538_not
g1195 not n540 ; n540_not
g1196 not a[20] ; a[20]_not
g1197 not b[20] ; b[20]_not
g1198 not n542 ; n542_not
g1199 not n543 ; n543_not
g1200 not n544 ; n544_not
g1201 not n541 ; n541_not
g1202 not n545 ; n545_not
g1203 not n546 ; n546_not
g1204 not n548 ; n548_not
g1205 not a[21] ; a[21]_not
g1206 not b[21] ; b[21]_not
g1207 not n550 ; n550_not
g1208 not n551 ; n551_not
g1209 not n552 ; n552_not
g1210 not n549 ; n549_not
g1211 not n553 ; n553_not
g1212 not n554 ; n554_not
g1213 not n556 ; n556_not
g1214 not a[22] ; a[22]_not
g1215 not b[22] ; b[22]_not
g1216 not n558 ; n558_not
g1217 not n559 ; n559_not
g1218 not n560 ; n560_not
g1219 not n557 ; n557_not
g1220 not n561 ; n561_not
g1221 not n562 ; n562_not
g1222 not n564 ; n564_not
g1223 not a[23] ; a[23]_not
g1224 not b[23] ; b[23]_not
g1225 not n566 ; n566_not
g1226 not n567 ; n567_not
g1227 not n568 ; n568_not
g1228 not n565 ; n565_not
g1229 not n569 ; n569_not
g1230 not n570 ; n570_not
g1231 not n572 ; n572_not
g1232 not a[24] ; a[24]_not
g1233 not b[24] ; b[24]_not
g1234 not n574 ; n574_not
g1235 not n575 ; n575_not
g1236 not n576 ; n576_not
g1237 not n573 ; n573_not
g1238 not n577 ; n577_not
g1239 not n578 ; n578_not
g1240 not n580 ; n580_not
g1241 not a[25] ; a[25]_not
g1242 not b[25] ; b[25]_not
g1243 not n582 ; n582_not
g1244 not n583 ; n583_not
g1245 not n584 ; n584_not
g1246 not n581 ; n581_not
g1247 not n585 ; n585_not
g1248 not n586 ; n586_not
g1249 not n588 ; n588_not
g1250 not a[26] ; a[26]_not
g1251 not b[26] ; b[26]_not
g1252 not n590 ; n590_not
g1253 not n591 ; n591_not
g1254 not n592 ; n592_not
g1255 not n589 ; n589_not
g1256 not n593 ; n593_not
g1257 not n594 ; n594_not
g1258 not n596 ; n596_not
g1259 not a[27] ; a[27]_not
g1260 not b[27] ; b[27]_not
g1261 not n598 ; n598_not
g1262 not n599 ; n599_not
g1263 not n600 ; n600_not
g1264 not n597 ; n597_not
g1265 not n601 ; n601_not
g1266 not n602 ; n602_not
g1267 not n604 ; n604_not
g1268 not a[28] ; a[28]_not
g1269 not b[28] ; b[28]_not
g1270 not n606 ; n606_not
g1271 not n607 ; n607_not
g1272 not n608 ; n608_not
g1273 not n605 ; n605_not
g1274 not n609 ; n609_not
g1275 not n610 ; n610_not
g1276 not n612 ; n612_not
g1277 not a[29] ; a[29]_not
g1278 not b[29] ; b[29]_not
g1279 not n614 ; n614_not
g1280 not n615 ; n615_not
g1281 not n616 ; n616_not
g1282 not n613 ; n613_not
g1283 not n617 ; n617_not
g1284 not n618 ; n618_not
g1285 not n620 ; n620_not
g1286 not a[30] ; a[30]_not
g1287 not b[30] ; b[30]_not
g1288 not n622 ; n622_not
g1289 not n623 ; n623_not
g1290 not n624 ; n624_not
g1291 not n621 ; n621_not
g1292 not n625 ; n625_not
g1293 not n626 ; n626_not
g1294 not n628 ; n628_not
g1295 not a[31] ; a[31]_not
g1296 not b[31] ; b[31]_not
g1297 not n630 ; n630_not
g1298 not n631 ; n631_not
g1299 not n632 ; n632_not
g1300 not n629 ; n629_not
g1301 not n633 ; n633_not
g1302 not n634 ; n634_not
g1303 not n636 ; n636_not
g1304 not a[32] ; a[32]_not
g1305 not b[32] ; b[32]_not
g1306 not n638 ; n638_not
g1307 not n639 ; n639_not
g1308 not n640 ; n640_not
g1309 not n637 ; n637_not
g1310 not n641 ; n641_not
g1311 not n642 ; n642_not
g1312 not n644 ; n644_not
g1313 not a[33] ; a[33]_not
g1314 not b[33] ; b[33]_not
g1315 not n646 ; n646_not
g1316 not n647 ; n647_not
g1317 not n648 ; n648_not
g1318 not n645 ; n645_not
g1319 not n649 ; n649_not
g1320 not n650 ; n650_not
g1321 not n652 ; n652_not
g1322 not a[34] ; a[34]_not
g1323 not b[34] ; b[34]_not
g1324 not n654 ; n654_not
g1325 not n655 ; n655_not
g1326 not n656 ; n656_not
g1327 not n653 ; n653_not
g1328 not n657 ; n657_not
g1329 not n658 ; n658_not
g1330 not n660 ; n660_not
g1331 not a[35] ; a[35]_not
g1332 not b[35] ; b[35]_not
g1333 not n662 ; n662_not
g1334 not n663 ; n663_not
g1335 not n664 ; n664_not
g1336 not n661 ; n661_not
g1337 not n665 ; n665_not
g1338 not n666 ; n666_not
g1339 not n668 ; n668_not
g1340 not a[36] ; a[36]_not
g1341 not b[36] ; b[36]_not
g1342 not n670 ; n670_not
g1343 not n671 ; n671_not
g1344 not n672 ; n672_not
g1345 not n669 ; n669_not
g1346 not n673 ; n673_not
g1347 not n674 ; n674_not
g1348 not n676 ; n676_not
g1349 not a[37] ; a[37]_not
g1350 not b[37] ; b[37]_not
g1351 not n678 ; n678_not
g1352 not n679 ; n679_not
g1353 not n680 ; n680_not
g1354 not n677 ; n677_not
g1355 not n681 ; n681_not
g1356 not n682 ; n682_not
g1357 not n684 ; n684_not
g1358 not a[38] ; a[38]_not
g1359 not b[38] ; b[38]_not
g1360 not n686 ; n686_not
g1361 not n687 ; n687_not
g1362 not n688 ; n688_not
g1363 not n685 ; n685_not
g1364 not n689 ; n689_not
g1365 not n690 ; n690_not
g1366 not n692 ; n692_not
g1367 not a[39] ; a[39]_not
g1368 not b[39] ; b[39]_not
g1369 not n694 ; n694_not
g1370 not n695 ; n695_not
g1371 not n696 ; n696_not
g1372 not n693 ; n693_not
g1373 not n697 ; n697_not
g1374 not n698 ; n698_not
g1375 not n700 ; n700_not
g1376 not a[40] ; a[40]_not
g1377 not b[40] ; b[40]_not
g1378 not n702 ; n702_not
g1379 not n703 ; n703_not
g1380 not n704 ; n704_not
g1381 not n701 ; n701_not
g1382 not n705 ; n705_not
g1383 not n706 ; n706_not
g1384 not n708 ; n708_not
g1385 not a[41] ; a[41]_not
g1386 not b[41] ; b[41]_not
g1387 not n710 ; n710_not
g1388 not n711 ; n711_not
g1389 not n712 ; n712_not
g1390 not n709 ; n709_not
g1391 not n713 ; n713_not
g1392 not n714 ; n714_not
g1393 not n716 ; n716_not
g1394 not a[42] ; a[42]_not
g1395 not b[42] ; b[42]_not
g1396 not n718 ; n718_not
g1397 not n719 ; n719_not
g1398 not n720 ; n720_not
g1399 not n717 ; n717_not
g1400 not n721 ; n721_not
g1401 not n722 ; n722_not
g1402 not n724 ; n724_not
g1403 not a[43] ; a[43]_not
g1404 not b[43] ; b[43]_not
g1405 not n726 ; n726_not
g1406 not n727 ; n727_not
g1407 not n728 ; n728_not
g1408 not n725 ; n725_not
g1409 not n729 ; n729_not
g1410 not n730 ; n730_not
g1411 not n732 ; n732_not
g1412 not a[44] ; a[44]_not
g1413 not b[44] ; b[44]_not
g1414 not n734 ; n734_not
g1415 not n735 ; n735_not
g1416 not n736 ; n736_not
g1417 not n733 ; n733_not
g1418 not n737 ; n737_not
g1419 not n738 ; n738_not
g1420 not n740 ; n740_not
g1421 not a[45] ; a[45]_not
g1422 not b[45] ; b[45]_not
g1423 not n742 ; n742_not
g1424 not n743 ; n743_not
g1425 not n744 ; n744_not
g1426 not n741 ; n741_not
g1427 not n745 ; n745_not
g1428 not n746 ; n746_not
g1429 not n748 ; n748_not
g1430 not a[46] ; a[46]_not
g1431 not b[46] ; b[46]_not
g1432 not n750 ; n750_not
g1433 not n751 ; n751_not
g1434 not n752 ; n752_not
g1435 not n749 ; n749_not
g1436 not n753 ; n753_not
g1437 not n754 ; n754_not
g1438 not n756 ; n756_not
g1439 not a[47] ; a[47]_not
g1440 not b[47] ; b[47]_not
g1441 not n758 ; n758_not
g1442 not n759 ; n759_not
g1443 not n760 ; n760_not
g1444 not n757 ; n757_not
g1445 not n761 ; n761_not
g1446 not n762 ; n762_not
g1447 not n764 ; n764_not
g1448 not a[48] ; a[48]_not
g1449 not b[48] ; b[48]_not
g1450 not n766 ; n766_not
g1451 not n767 ; n767_not
g1452 not n768 ; n768_not
g1453 not n765 ; n765_not
g1454 not n769 ; n769_not
g1455 not n770 ; n770_not
g1456 not n772 ; n772_not
g1457 not a[49] ; a[49]_not
g1458 not b[49] ; b[49]_not
g1459 not n774 ; n774_not
g1460 not n775 ; n775_not
g1461 not n776 ; n776_not
g1462 not n773 ; n773_not
g1463 not n777 ; n777_not
g1464 not n778 ; n778_not
g1465 not n780 ; n780_not
g1466 not a[50] ; a[50]_not
g1467 not b[50] ; b[50]_not
g1468 not n782 ; n782_not
g1469 not n783 ; n783_not
g1470 not n784 ; n784_not
g1471 not n781 ; n781_not
g1472 not n785 ; n785_not
g1473 not n786 ; n786_not
g1474 not n788 ; n788_not
g1475 not a[51] ; a[51]_not
g1476 not b[51] ; b[51]_not
g1477 not n790 ; n790_not
g1478 not n791 ; n791_not
g1479 not n792 ; n792_not
g1480 not n789 ; n789_not
g1481 not n793 ; n793_not
g1482 not n794 ; n794_not
g1483 not n796 ; n796_not
g1484 not a[52] ; a[52]_not
g1485 not b[52] ; b[52]_not
g1486 not n798 ; n798_not
g1487 not n799 ; n799_not
g1488 not n800 ; n800_not
g1489 not n797 ; n797_not
g1490 not n801 ; n801_not
g1491 not n802 ; n802_not
g1492 not n804 ; n804_not
g1493 not a[53] ; a[53]_not
g1494 not b[53] ; b[53]_not
g1495 not n806 ; n806_not
g1496 not n807 ; n807_not
g1497 not n808 ; n808_not
g1498 not n805 ; n805_not
g1499 not n809 ; n809_not
g1500 not n810 ; n810_not
g1501 not n812 ; n812_not
g1502 not a[54] ; a[54]_not
g1503 not b[54] ; b[54]_not
g1504 not n814 ; n814_not
g1505 not n815 ; n815_not
g1506 not n816 ; n816_not
g1507 not n813 ; n813_not
g1508 not n817 ; n817_not
g1509 not n818 ; n818_not
g1510 not n820 ; n820_not
g1511 not a[55] ; a[55]_not
g1512 not b[55] ; b[55]_not
g1513 not n822 ; n822_not
g1514 not n823 ; n823_not
g1515 not n824 ; n824_not
g1516 not n821 ; n821_not
g1517 not n825 ; n825_not
g1518 not n826 ; n826_not
g1519 not n828 ; n828_not
g1520 not a[56] ; a[56]_not
g1521 not b[56] ; b[56]_not
g1522 not n830 ; n830_not
g1523 not n831 ; n831_not
g1524 not n832 ; n832_not
g1525 not n829 ; n829_not
g1526 not n833 ; n833_not
g1527 not n834 ; n834_not
g1528 not n836 ; n836_not
g1529 not a[57] ; a[57]_not
g1530 not b[57] ; b[57]_not
g1531 not n838 ; n838_not
g1532 not n839 ; n839_not
g1533 not n840 ; n840_not
g1534 not n837 ; n837_not
g1535 not n841 ; n841_not
g1536 not n842 ; n842_not
g1537 not n844 ; n844_not
g1538 not a[58] ; a[58]_not
g1539 not b[58] ; b[58]_not
g1540 not n846 ; n846_not
g1541 not n847 ; n847_not
g1542 not n848 ; n848_not
g1543 not n845 ; n845_not
g1544 not n849 ; n849_not
g1545 not n850 ; n850_not
g1546 not n852 ; n852_not
g1547 not a[59] ; a[59]_not
g1548 not b[59] ; b[59]_not
g1549 not n854 ; n854_not
g1550 not n855 ; n855_not
g1551 not n856 ; n856_not
g1552 not n853 ; n853_not
g1553 not n857 ; n857_not
g1554 not n858 ; n858_not
g1555 not n860 ; n860_not
g1556 not a[60] ; a[60]_not
g1557 not b[60] ; b[60]_not
g1558 not n862 ; n862_not
g1559 not n863 ; n863_not
g1560 not n864 ; n864_not
g1561 not n861 ; n861_not
g1562 not n865 ; n865_not
g1563 not n866 ; n866_not
g1564 not n868 ; n868_not
g1565 not a[61] ; a[61]_not
g1566 not b[61] ; b[61]_not
g1567 not n870 ; n870_not
g1568 not n871 ; n871_not
g1569 not n872 ; n872_not
g1570 not n869 ; n869_not
g1571 not n873 ; n873_not
g1572 not n874 ; n874_not
g1573 not n876 ; n876_not
g1574 not a[62] ; a[62]_not
g1575 not b[62] ; b[62]_not
g1576 not n878 ; n878_not
g1577 not n879 ; n879_not
g1578 not n880 ; n880_not
g1579 not n877 ; n877_not
g1580 not n881 ; n881_not
g1581 not n882 ; n882_not
g1582 not n884 ; n884_not
g1583 not a[63] ; a[63]_not
g1584 not b[63] ; b[63]_not
g1585 not n886 ; n886_not
g1586 not n887 ; n887_not
g1587 not n888 ; n888_not
g1588 not n885 ; n885_not
g1589 not n889 ; n889_not
g1590 not n890 ; n890_not
g1591 not n892 ; n892_not
g1592 not a[64] ; a[64]_not
g1593 not b[64] ; b[64]_not
g1594 not n894 ; n894_not
g1595 not n895 ; n895_not
g1596 not n896 ; n896_not
g1597 not n893 ; n893_not
g1598 not n897 ; n897_not
g1599 not n898 ; n898_not
g1600 not n900 ; n900_not
g1601 not a[65] ; a[65]_not
g1602 not b[65] ; b[65]_not
g1603 not n902 ; n902_not
g1604 not n903 ; n903_not
g1605 not n904 ; n904_not
g1606 not n901 ; n901_not
g1607 not n905 ; n905_not
g1608 not n906 ; n906_not
g1609 not n908 ; n908_not
g1610 not a[66] ; a[66]_not
g1611 not b[66] ; b[66]_not
g1612 not n910 ; n910_not
g1613 not n911 ; n911_not
g1614 not n912 ; n912_not
g1615 not n909 ; n909_not
g1616 not n913 ; n913_not
g1617 not n914 ; n914_not
g1618 not n916 ; n916_not
g1619 not a[67] ; a[67]_not
g1620 not b[67] ; b[67]_not
g1621 not n918 ; n918_not
g1622 not n919 ; n919_not
g1623 not n920 ; n920_not
g1624 not n917 ; n917_not
g1625 not n921 ; n921_not
g1626 not n922 ; n922_not
g1627 not n924 ; n924_not
g1628 not a[68] ; a[68]_not
g1629 not b[68] ; b[68]_not
g1630 not n926 ; n926_not
g1631 not n927 ; n927_not
g1632 not n928 ; n928_not
g1633 not n925 ; n925_not
g1634 not n929 ; n929_not
g1635 not n930 ; n930_not
g1636 not n932 ; n932_not
g1637 not a[69] ; a[69]_not
g1638 not b[69] ; b[69]_not
g1639 not n934 ; n934_not
g1640 not n935 ; n935_not
g1641 not n936 ; n936_not
g1642 not n933 ; n933_not
g1643 not n937 ; n937_not
g1644 not n938 ; n938_not
g1645 not n940 ; n940_not
g1646 not a[70] ; a[70]_not
g1647 not b[70] ; b[70]_not
g1648 not n942 ; n942_not
g1649 not n943 ; n943_not
g1650 not n944 ; n944_not
g1651 not n941 ; n941_not
g1652 not n945 ; n945_not
g1653 not n946 ; n946_not
g1654 not n948 ; n948_not
g1655 not a[71] ; a[71]_not
g1656 not b[71] ; b[71]_not
g1657 not n950 ; n950_not
g1658 not n951 ; n951_not
g1659 not n952 ; n952_not
g1660 not n949 ; n949_not
g1661 not n953 ; n953_not
g1662 not n954 ; n954_not
g1663 not n956 ; n956_not
g1664 not a[72] ; a[72]_not
g1665 not b[72] ; b[72]_not
g1666 not n958 ; n958_not
g1667 not n959 ; n959_not
g1668 not n960 ; n960_not
g1669 not n957 ; n957_not
g1670 not n961 ; n961_not
g1671 not n962 ; n962_not
g1672 not n964 ; n964_not
g1673 not a[73] ; a[73]_not
g1674 not b[73] ; b[73]_not
g1675 not n966 ; n966_not
g1676 not n967 ; n967_not
g1677 not n968 ; n968_not
g1678 not n965 ; n965_not
g1679 not n969 ; n969_not
g1680 not n970 ; n970_not
g1681 not n972 ; n972_not
g1682 not a[74] ; a[74]_not
g1683 not b[74] ; b[74]_not
g1684 not n974 ; n974_not
g1685 not n975 ; n975_not
g1686 not n976 ; n976_not
g1687 not n973 ; n973_not
g1688 not n977 ; n977_not
g1689 not n978 ; n978_not
g1690 not n980 ; n980_not
g1691 not a[75] ; a[75]_not
g1692 not b[75] ; b[75]_not
g1693 not n982 ; n982_not
g1694 not n983 ; n983_not
g1695 not n984 ; n984_not
g1696 not n981 ; n981_not
g1697 not n985 ; n985_not
g1698 not n986 ; n986_not
g1699 not n988 ; n988_not
g1700 not a[76] ; a[76]_not
g1701 not b[76] ; b[76]_not
g1702 not n990 ; n990_not
g1703 not n991 ; n991_not
g1704 not n992 ; n992_not
g1705 not n989 ; n989_not
g1706 not n993 ; n993_not
g1707 not n994 ; n994_not
g1708 not n996 ; n996_not
g1709 not a[77] ; a[77]_not
g1710 not b[77] ; b[77]_not
g1711 not n998 ; n998_not
g1712 not n999 ; n999_not
g1713 not n1000 ; n1000_not
g1714 not n997 ; n997_not
g1715 not n1001 ; n1001_not
g1716 not n1002 ; n1002_not
g1717 not n1004 ; n1004_not
g1718 not a[78] ; a[78]_not
g1719 not b[78] ; b[78]_not
g1720 not n1006 ; n1006_not
g1721 not n1007 ; n1007_not
g1722 not n1008 ; n1008_not
g1723 not n1005 ; n1005_not
g1724 not n1009 ; n1009_not
g1725 not n1010 ; n1010_not
g1726 not n1012 ; n1012_not
g1727 not a[79] ; a[79]_not
g1728 not b[79] ; b[79]_not
g1729 not n1014 ; n1014_not
g1730 not n1015 ; n1015_not
g1731 not n1016 ; n1016_not
g1732 not n1013 ; n1013_not
g1733 not n1017 ; n1017_not
g1734 not n1018 ; n1018_not
g1735 not n1020 ; n1020_not
g1736 not a[80] ; a[80]_not
g1737 not b[80] ; b[80]_not
g1738 not n1022 ; n1022_not
g1739 not n1023 ; n1023_not
g1740 not n1024 ; n1024_not
g1741 not n1021 ; n1021_not
g1742 not n1025 ; n1025_not
g1743 not n1026 ; n1026_not
g1744 not n1028 ; n1028_not
g1745 not a[81] ; a[81]_not
g1746 not b[81] ; b[81]_not
g1747 not n1030 ; n1030_not
g1748 not n1031 ; n1031_not
g1749 not n1032 ; n1032_not
g1750 not n1029 ; n1029_not
g1751 not n1033 ; n1033_not
g1752 not n1034 ; n1034_not
g1753 not n1036 ; n1036_not
g1754 not a[82] ; a[82]_not
g1755 not b[82] ; b[82]_not
g1756 not n1038 ; n1038_not
g1757 not n1039 ; n1039_not
g1758 not n1040 ; n1040_not
g1759 not n1037 ; n1037_not
g1760 not n1041 ; n1041_not
g1761 not n1042 ; n1042_not
g1762 not n1044 ; n1044_not
g1763 not a[83] ; a[83]_not
g1764 not b[83] ; b[83]_not
g1765 not n1046 ; n1046_not
g1766 not n1047 ; n1047_not
g1767 not n1048 ; n1048_not
g1768 not n1045 ; n1045_not
g1769 not n1049 ; n1049_not
g1770 not n1050 ; n1050_not
g1771 not n1052 ; n1052_not
g1772 not a[84] ; a[84]_not
g1773 not b[84] ; b[84]_not
g1774 not n1054 ; n1054_not
g1775 not n1055 ; n1055_not
g1776 not n1056 ; n1056_not
g1777 not n1053 ; n1053_not
g1778 not n1057 ; n1057_not
g1779 not n1058 ; n1058_not
g1780 not n1060 ; n1060_not
g1781 not a[85] ; a[85]_not
g1782 not b[85] ; b[85]_not
g1783 not n1062 ; n1062_not
g1784 not n1063 ; n1063_not
g1785 not n1064 ; n1064_not
g1786 not n1061 ; n1061_not
g1787 not n1065 ; n1065_not
g1788 not n1066 ; n1066_not
g1789 not n1068 ; n1068_not
g1790 not a[86] ; a[86]_not
g1791 not b[86] ; b[86]_not
g1792 not n1070 ; n1070_not
g1793 not n1071 ; n1071_not
g1794 not n1072 ; n1072_not
g1795 not n1069 ; n1069_not
g1796 not n1073 ; n1073_not
g1797 not n1074 ; n1074_not
g1798 not n1076 ; n1076_not
g1799 not a[87] ; a[87]_not
g1800 not b[87] ; b[87]_not
g1801 not n1078 ; n1078_not
g1802 not n1079 ; n1079_not
g1803 not n1080 ; n1080_not
g1804 not n1077 ; n1077_not
g1805 not n1081 ; n1081_not
g1806 not n1082 ; n1082_not
g1807 not n1084 ; n1084_not
g1808 not a[88] ; a[88]_not
g1809 not b[88] ; b[88]_not
g1810 not n1086 ; n1086_not
g1811 not n1087 ; n1087_not
g1812 not n1088 ; n1088_not
g1813 not n1085 ; n1085_not
g1814 not n1089 ; n1089_not
g1815 not n1090 ; n1090_not
g1816 not n1092 ; n1092_not
g1817 not a[89] ; a[89]_not
g1818 not b[89] ; b[89]_not
g1819 not n1094 ; n1094_not
g1820 not n1095 ; n1095_not
g1821 not n1096 ; n1096_not
g1822 not n1093 ; n1093_not
g1823 not n1097 ; n1097_not
g1824 not n1098 ; n1098_not
g1825 not n1100 ; n1100_not
g1826 not a[90] ; a[90]_not
g1827 not b[90] ; b[90]_not
g1828 not n1102 ; n1102_not
g1829 not n1103 ; n1103_not
g1830 not n1104 ; n1104_not
g1831 not n1101 ; n1101_not
g1832 not n1105 ; n1105_not
g1833 not n1106 ; n1106_not
g1834 not n1108 ; n1108_not
g1835 not a[91] ; a[91]_not
g1836 not b[91] ; b[91]_not
g1837 not n1110 ; n1110_not
g1838 not n1111 ; n1111_not
g1839 not n1112 ; n1112_not
g1840 not n1109 ; n1109_not
g1841 not n1113 ; n1113_not
g1842 not n1114 ; n1114_not
g1843 not n1116 ; n1116_not
g1844 not a[92] ; a[92]_not
g1845 not b[92] ; b[92]_not
g1846 not n1118 ; n1118_not
g1847 not n1119 ; n1119_not
g1848 not n1120 ; n1120_not
g1849 not n1117 ; n1117_not
g1850 not n1121 ; n1121_not
g1851 not n1122 ; n1122_not
g1852 not n1124 ; n1124_not
g1853 not a[93] ; a[93]_not
g1854 not b[93] ; b[93]_not
g1855 not n1126 ; n1126_not
g1856 not n1127 ; n1127_not
g1857 not n1128 ; n1128_not
g1858 not n1125 ; n1125_not
g1859 not n1129 ; n1129_not
g1860 not n1130 ; n1130_not
g1861 not n1132 ; n1132_not
g1862 not a[94] ; a[94]_not
g1863 not b[94] ; b[94]_not
g1864 not n1134 ; n1134_not
g1865 not n1135 ; n1135_not
g1866 not n1136 ; n1136_not
g1867 not n1133 ; n1133_not
g1868 not n1137 ; n1137_not
g1869 not n1138 ; n1138_not
g1870 not n1140 ; n1140_not
g1871 not a[95] ; a[95]_not
g1872 not b[95] ; b[95]_not
g1873 not n1142 ; n1142_not
g1874 not n1143 ; n1143_not
g1875 not n1144 ; n1144_not
g1876 not n1141 ; n1141_not
g1877 not n1145 ; n1145_not
g1878 not n1146 ; n1146_not
g1879 not n1148 ; n1148_not
g1880 not a[96] ; a[96]_not
g1881 not b[96] ; b[96]_not
g1882 not n1150 ; n1150_not
g1883 not n1151 ; n1151_not
g1884 not n1152 ; n1152_not
g1885 not n1149 ; n1149_not
g1886 not n1153 ; n1153_not
g1887 not n1154 ; n1154_not
g1888 not n1156 ; n1156_not
g1889 not a[97] ; a[97]_not
g1890 not b[97] ; b[97]_not
g1891 not n1158 ; n1158_not
g1892 not n1159 ; n1159_not
g1893 not n1160 ; n1160_not
g1894 not n1157 ; n1157_not
g1895 not n1161 ; n1161_not
g1896 not n1162 ; n1162_not
g1897 not n1164 ; n1164_not
g1898 not a[98] ; a[98]_not
g1899 not b[98] ; b[98]_not
g1900 not n1166 ; n1166_not
g1901 not n1167 ; n1167_not
g1902 not n1168 ; n1168_not
g1903 not n1165 ; n1165_not
g1904 not n1169 ; n1169_not
g1905 not n1170 ; n1170_not
g1906 not n1172 ; n1172_not
g1907 not a[99] ; a[99]_not
g1908 not b[99] ; b[99]_not
g1909 not n1174 ; n1174_not
g1910 not n1175 ; n1175_not
g1911 not n1176 ; n1176_not
g1912 not n1173 ; n1173_not
g1913 not n1177 ; n1177_not
g1914 not n1178 ; n1178_not
g1915 not n1180 ; n1180_not
g1916 not a[100] ; a[100]_not
g1917 not b[100] ; b[100]_not
g1918 not n1182 ; n1182_not
g1919 not n1183 ; n1183_not
g1920 not n1184 ; n1184_not
g1921 not n1181 ; n1181_not
g1922 not n1185 ; n1185_not
g1923 not n1186 ; n1186_not
g1924 not n1188 ; n1188_not
g1925 not a[101] ; a[101]_not
g1926 not b[101] ; b[101]_not
g1927 not n1190 ; n1190_not
g1928 not n1191 ; n1191_not
g1929 not n1192 ; n1192_not
g1930 not n1189 ; n1189_not
g1931 not n1193 ; n1193_not
g1932 not n1194 ; n1194_not
g1933 not n1196 ; n1196_not
g1934 not a[102] ; a[102]_not
g1935 not b[102] ; b[102]_not
g1936 not n1198 ; n1198_not
g1937 not n1199 ; n1199_not
g1938 not n1200 ; n1200_not
g1939 not n1197 ; n1197_not
g1940 not n1201 ; n1201_not
g1941 not n1202 ; n1202_not
g1942 not n1204 ; n1204_not
g1943 not a[103] ; a[103]_not
g1944 not b[103] ; b[103]_not
g1945 not n1206 ; n1206_not
g1946 not n1207 ; n1207_not
g1947 not n1208 ; n1208_not
g1948 not n1205 ; n1205_not
g1949 not n1209 ; n1209_not
g1950 not n1210 ; n1210_not
g1951 not n1212 ; n1212_not
g1952 not a[104] ; a[104]_not
g1953 not b[104] ; b[104]_not
g1954 not n1214 ; n1214_not
g1955 not n1215 ; n1215_not
g1956 not n1216 ; n1216_not
g1957 not n1213 ; n1213_not
g1958 not n1217 ; n1217_not
g1959 not n1218 ; n1218_not
g1960 not n1220 ; n1220_not
g1961 not a[105] ; a[105]_not
g1962 not b[105] ; b[105]_not
g1963 not n1222 ; n1222_not
g1964 not n1223 ; n1223_not
g1965 not n1224 ; n1224_not
g1966 not n1221 ; n1221_not
g1967 not n1225 ; n1225_not
g1968 not n1226 ; n1226_not
g1969 not n1228 ; n1228_not
g1970 not a[106] ; a[106]_not
g1971 not b[106] ; b[106]_not
g1972 not n1230 ; n1230_not
g1973 not n1231 ; n1231_not
g1974 not n1232 ; n1232_not
g1975 not n1229 ; n1229_not
g1976 not n1233 ; n1233_not
g1977 not n1234 ; n1234_not
g1978 not n1236 ; n1236_not
g1979 not a[107] ; a[107]_not
g1980 not b[107] ; b[107]_not
g1981 not n1238 ; n1238_not
g1982 not n1239 ; n1239_not
g1983 not n1240 ; n1240_not
g1984 not n1237 ; n1237_not
g1985 not n1241 ; n1241_not
g1986 not n1242 ; n1242_not
g1987 not n1244 ; n1244_not
g1988 not a[108] ; a[108]_not
g1989 not b[108] ; b[108]_not
g1990 not n1246 ; n1246_not
g1991 not n1247 ; n1247_not
g1992 not n1248 ; n1248_not
g1993 not n1245 ; n1245_not
g1994 not n1249 ; n1249_not
g1995 not n1250 ; n1250_not
g1996 not n1252 ; n1252_not
g1997 not a[109] ; a[109]_not
g1998 not b[109] ; b[109]_not
g1999 not n1254 ; n1254_not
g2000 not n1255 ; n1255_not
g2001 not n1256 ; n1256_not
g2002 not n1253 ; n1253_not
g2003 not n1257 ; n1257_not
g2004 not n1258 ; n1258_not
g2005 not n1260 ; n1260_not
g2006 not a[110] ; a[110]_not
g2007 not b[110] ; b[110]_not
g2008 not n1262 ; n1262_not
g2009 not n1263 ; n1263_not
g2010 not n1264 ; n1264_not
g2011 not n1261 ; n1261_not
g2012 not n1265 ; n1265_not
g2013 not n1266 ; n1266_not
g2014 not n1268 ; n1268_not
g2015 not a[111] ; a[111]_not
g2016 not b[111] ; b[111]_not
g2017 not n1270 ; n1270_not
g2018 not n1271 ; n1271_not
g2019 not n1272 ; n1272_not
g2020 not n1269 ; n1269_not
g2021 not n1273 ; n1273_not
g2022 not n1274 ; n1274_not
g2023 not n1276 ; n1276_not
g2024 not a[112] ; a[112]_not
g2025 not b[112] ; b[112]_not
g2026 not n1278 ; n1278_not
g2027 not n1279 ; n1279_not
g2028 not n1280 ; n1280_not
g2029 not n1277 ; n1277_not
g2030 not n1281 ; n1281_not
g2031 not n1282 ; n1282_not
g2032 not n1284 ; n1284_not
g2033 not a[113] ; a[113]_not
g2034 not b[113] ; b[113]_not
g2035 not n1286 ; n1286_not
g2036 not n1287 ; n1287_not
g2037 not n1288 ; n1288_not
g2038 not n1285 ; n1285_not
g2039 not n1289 ; n1289_not
g2040 not n1290 ; n1290_not
g2041 not n1292 ; n1292_not
g2042 not a[114] ; a[114]_not
g2043 not b[114] ; b[114]_not
g2044 not n1294 ; n1294_not
g2045 not n1295 ; n1295_not
g2046 not n1296 ; n1296_not
g2047 not n1293 ; n1293_not
g2048 not n1297 ; n1297_not
g2049 not n1298 ; n1298_not
g2050 not n1300 ; n1300_not
g2051 not a[115] ; a[115]_not
g2052 not b[115] ; b[115]_not
g2053 not n1302 ; n1302_not
g2054 not n1303 ; n1303_not
g2055 not n1304 ; n1304_not
g2056 not n1301 ; n1301_not
g2057 not n1305 ; n1305_not
g2058 not n1306 ; n1306_not
g2059 not n1308 ; n1308_not
g2060 not a[116] ; a[116]_not
g2061 not b[116] ; b[116]_not
g2062 not n1310 ; n1310_not
g2063 not n1311 ; n1311_not
g2064 not n1312 ; n1312_not
g2065 not n1309 ; n1309_not
g2066 not n1313 ; n1313_not
g2067 not n1314 ; n1314_not
g2068 not n1316 ; n1316_not
g2069 not a[117] ; a[117]_not
g2070 not b[117] ; b[117]_not
g2071 not n1318 ; n1318_not
g2072 not n1319 ; n1319_not
g2073 not n1320 ; n1320_not
g2074 not n1317 ; n1317_not
g2075 not n1321 ; n1321_not
g2076 not n1322 ; n1322_not
g2077 not n1324 ; n1324_not
g2078 not a[118] ; a[118]_not
g2079 not b[118] ; b[118]_not
g2080 not n1326 ; n1326_not
g2081 not n1327 ; n1327_not
g2082 not n1328 ; n1328_not
g2083 not n1325 ; n1325_not
g2084 not n1329 ; n1329_not
g2085 not n1330 ; n1330_not
g2086 not n1332 ; n1332_not
g2087 not a[119] ; a[119]_not
g2088 not b[119] ; b[119]_not
g2089 not n1334 ; n1334_not
g2090 not n1335 ; n1335_not
g2091 not n1336 ; n1336_not
g2092 not n1333 ; n1333_not
g2093 not n1337 ; n1337_not
g2094 not n1338 ; n1338_not
g2095 not n1340 ; n1340_not
g2096 not a[120] ; a[120]_not
g2097 not b[120] ; b[120]_not
g2098 not n1342 ; n1342_not
g2099 not n1343 ; n1343_not
g2100 not n1344 ; n1344_not
g2101 not n1341 ; n1341_not
g2102 not n1345 ; n1345_not
g2103 not n1346 ; n1346_not
g2104 not n1348 ; n1348_not
g2105 not a[121] ; a[121]_not
g2106 not b[121] ; b[121]_not
g2107 not n1350 ; n1350_not
g2108 not n1351 ; n1351_not
g2109 not n1352 ; n1352_not
g2110 not n1349 ; n1349_not
g2111 not n1353 ; n1353_not
g2112 not n1354 ; n1354_not
g2113 not n1356 ; n1356_not
g2114 not a[122] ; a[122]_not
g2115 not b[122] ; b[122]_not
g2116 not n1358 ; n1358_not
g2117 not n1359 ; n1359_not
g2118 not n1360 ; n1360_not
g2119 not n1357 ; n1357_not
g2120 not n1361 ; n1361_not
g2121 not n1362 ; n1362_not
g2122 not n1364 ; n1364_not
g2123 not a[123] ; a[123]_not
g2124 not b[123] ; b[123]_not
g2125 not n1366 ; n1366_not
g2126 not n1367 ; n1367_not
g2127 not n1368 ; n1368_not
g2128 not n1365 ; n1365_not
g2129 not n1369 ; n1369_not
g2130 not n1370 ; n1370_not
g2131 not n1372 ; n1372_not
g2132 not a[124] ; a[124]_not
g2133 not b[124] ; b[124]_not
g2134 not n1374 ; n1374_not
g2135 not n1375 ; n1375_not
g2136 not n1376 ; n1376_not
g2137 not n1373 ; n1373_not
g2138 not n1377 ; n1377_not
g2139 not n1378 ; n1378_not
g2140 not n1380 ; n1380_not
g2141 not a[125] ; a[125]_not
g2142 not b[125] ; b[125]_not
g2143 not n1382 ; n1382_not
g2144 not n1383 ; n1383_not
g2145 not n1384 ; n1384_not
g2146 not n1381 ; n1381_not
g2147 not n1385 ; n1385_not
g2148 not n1386 ; n1386_not
g2149 not n1388 ; n1388_not
g2150 not a[126] ; a[126]_not
g2151 not b[126] ; b[126]_not
g2152 not n1390 ; n1390_not
g2153 not n1391 ; n1391_not
g2154 not n1392 ; n1392_not
g2155 not n1389 ; n1389_not
g2156 not n1393 ; n1393_not
g2157 not n1394 ; n1394_not
g2158 not n1396 ; n1396_not
g2159 not a[127] ; a[127]_not
g2160 not b[127] ; b[127]_not
g2161 not n1398 ; n1398_not
g2162 not n1399 ; n1399_not
g2163 not n1400 ; n1400_not
g2164 not n1397 ; n1397_not
g2165 not n1401 ; n1401_not
g2166 not n1402 ; n1402_not
g2167 not n1404 ; n1404_not
o f[0]
o f[1]
o f[2]
o f[3]
o f[4]
o f[5]
o f[6]
o f[7]
o f[8]
o f[9]
o f[10]
o f[11]
o f[12]
o f[13]
o f[14]
o f[15]
o f[16]
o f[17]
o f[18]
o f[19]
o f[20]
o f[21]
o f[22]
o f[23]
o f[24]
o f[25]
o f[26]
o f[27]
o f[28]
o f[29]
o f[30]
o f[31]
o f[32]
o f[33]
o f[34]
o f[35]
o f[36]
o f[37]
o f[38]
o f[39]
o f[40]
o f[41]
o f[42]
o f[43]
o f[44]
o f[45]
o f[46]
o f[47]
o f[48]
o f[49]
o f[50]
o f[51]
o f[52]
o f[53]
o f[54]
o f[55]
o f[56]
o f[57]
o f[58]
o f[59]
o f[60]
o f[61]
o f[62]
o f[63]
o f[64]
o f[65]
o f[66]
o f[67]
o f[68]
o f[69]
o f[70]
o f[71]
o f[72]
o f[73]
o f[74]
o f[75]
o f[76]
o f[77]
o f[78]
o f[79]
o f[80]
o f[81]
o f[82]
o f[83]
o f[84]
o f[85]
o f[86]
o f[87]
o f[88]
o f[89]
o f[90]
o f[91]
o f[92]
o f[93]
o f[94]
o f[95]
o f[96]
o f[97]
o f[98]
o f[99]
o f[100]
o f[101]
o f[102]
o f[103]
o f[104]
o f[105]
o f[106]
o f[107]
o f[108]
o f[109]
o f[110]
o f[111]
o f[112]
o f[113]
o f[114]
o f[115]
o f[116]
o f[117]
o f[118]
o f[119]
o f[120]
o f[121]
o f[122]
o f[123]
o f[124]
o f[125]
o f[126]
o f[127]
o cOut
